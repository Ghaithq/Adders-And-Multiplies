
module register_N32_2 ( clk, reset, reg_in, reg_out );
  input [31:0] reg_in;
  output [31:0] reg_out;
  input clk, reset;
  wire   n33, n34, n35, n36;

  SDFF_X1 reg_out_reg_31_ ( .D(1'b0), .SI(n33), .SE(reg_in[31]), .CK(clk), .Q(
        reg_out[31]) );
  SDFF_X1 reg_out_reg_30_ ( .D(1'b0), .SI(n33), .SE(reg_in[30]), .CK(clk), .Q(
        reg_out[30]) );
  SDFF_X1 reg_out_reg_29_ ( .D(1'b0), .SI(n33), .SE(reg_in[29]), .CK(clk), .Q(
        reg_out[29]) );
  SDFF_X1 reg_out_reg_28_ ( .D(1'b0), .SI(n33), .SE(reg_in[28]), .CK(clk), .Q(
        reg_out[28]) );
  SDFF_X1 reg_out_reg_27_ ( .D(1'b0), .SI(n33), .SE(reg_in[27]), .CK(clk), .Q(
        reg_out[27]) );
  SDFF_X1 reg_out_reg_26_ ( .D(1'b0), .SI(n33), .SE(reg_in[26]), .CK(clk), .Q(
        reg_out[26]) );
  SDFF_X1 reg_out_reg_25_ ( .D(1'b0), .SI(n33), .SE(reg_in[25]), .CK(clk), .Q(
        reg_out[25]) );
  SDFF_X1 reg_out_reg_24_ ( .D(1'b0), .SI(n33), .SE(reg_in[24]), .CK(clk), .Q(
        reg_out[24]) );
  SDFF_X1 reg_out_reg_23_ ( .D(1'b0), .SI(n33), .SE(reg_in[23]), .CK(clk), .Q(
        reg_out[23]) );
  SDFF_X1 reg_out_reg_22_ ( .D(1'b0), .SI(n33), .SE(reg_in[22]), .CK(clk), .Q(
        reg_out[22]) );
  SDFF_X1 reg_out_reg_21_ ( .D(1'b0), .SI(n33), .SE(reg_in[21]), .CK(clk), .Q(
        reg_out[21]) );
  SDFF_X1 reg_out_reg_20_ ( .D(1'b0), .SI(n34), .SE(reg_in[20]), .CK(clk), .Q(
        reg_out[20]) );
  SDFF_X1 reg_out_reg_19_ ( .D(1'b0), .SI(n34), .SE(reg_in[19]), .CK(clk), .Q(
        reg_out[19]) );
  SDFF_X1 reg_out_reg_18_ ( .D(1'b0), .SI(n34), .SE(reg_in[18]), .CK(clk), .Q(
        reg_out[18]) );
  SDFF_X1 reg_out_reg_17_ ( .D(1'b0), .SI(n34), .SE(reg_in[17]), .CK(clk), .Q(
        reg_out[17]) );
  SDFF_X1 reg_out_reg_16_ ( .D(1'b0), .SI(n34), .SE(reg_in[16]), .CK(clk), .Q(
        reg_out[16]) );
  SDFF_X1 reg_out_reg_15_ ( .D(1'b0), .SI(n34), .SE(reg_in[15]), .CK(clk), .Q(
        reg_out[15]) );
  SDFF_X1 reg_out_reg_14_ ( .D(1'b0), .SI(n34), .SE(reg_in[14]), .CK(clk), .Q(
        reg_out[14]) );
  SDFF_X1 reg_out_reg_13_ ( .D(1'b0), .SI(n34), .SE(reg_in[13]), .CK(clk), .Q(
        reg_out[13]) );
  SDFF_X1 reg_out_reg_12_ ( .D(1'b0), .SI(n34), .SE(reg_in[12]), .CK(clk), .Q(
        reg_out[12]) );
  SDFF_X1 reg_out_reg_11_ ( .D(1'b0), .SI(n34), .SE(reg_in[11]), .CK(clk), .Q(
        reg_out[11]) );
  SDFF_X1 reg_out_reg_10_ ( .D(1'b0), .SI(n34), .SE(reg_in[10]), .CK(clk), .Q(
        reg_out[10]) );
  SDFF_X1 reg_out_reg_9_ ( .D(1'b0), .SI(n35), .SE(reg_in[9]), .CK(clk), .Q(
        reg_out[9]) );
  SDFF_X1 reg_out_reg_8_ ( .D(1'b0), .SI(n35), .SE(reg_in[8]), .CK(clk), .Q(
        reg_out[8]) );
  SDFF_X1 reg_out_reg_7_ ( .D(1'b0), .SI(n35), .SE(reg_in[7]), .CK(clk), .Q(
        reg_out[7]) );
  SDFF_X1 reg_out_reg_6_ ( .D(1'b0), .SI(n35), .SE(reg_in[6]), .CK(clk), .Q(
        reg_out[6]) );
  SDFF_X1 reg_out_reg_5_ ( .D(1'b0), .SI(n35), .SE(reg_in[5]), .CK(clk), .Q(
        reg_out[5]) );
  SDFF_X1 reg_out_reg_4_ ( .D(1'b0), .SI(n35), .SE(reg_in[4]), .CK(clk), .Q(
        reg_out[4]) );
  SDFF_X1 reg_out_reg_3_ ( .D(1'b0), .SI(n35), .SE(reg_in[3]), .CK(clk), .Q(
        reg_out[3]) );
  SDFF_X1 reg_out_reg_2_ ( .D(1'b0), .SI(n35), .SE(reg_in[2]), .CK(clk), .Q(
        reg_out[2]) );
  SDFF_X1 reg_out_reg_1_ ( .D(1'b0), .SI(n35), .SE(reg_in[1]), .CK(clk), .Q(
        reg_out[1]) );
  SDFF_X1 reg_out_reg_0_ ( .D(1'b0), .SI(n35), .SE(reg_in[0]), .CK(clk), .Q(
        reg_out[0]) );
  BUF_X1 U35 ( .A(n36), .Z(n34) );
  BUF_X1 U36 ( .A(n36), .Z(n33) );
  BUF_X1 U37 ( .A(n36), .Z(n35) );
  INV_X1 U38 ( .A(reset), .ZN(n36) );
endmodule


module register_N32_3 ( clk, reset, reg_in, reg_out );
  input [31:0] reg_in;
  output [31:0] reg_out;
  input clk, reset;
  wire   n33, n34, n35, n36;

  SDFF_X1 reg_out_reg_31_ ( .D(1'b0), .SI(n33), .SE(reg_in[31]), .CK(clk), .Q(
        reg_out[31]) );
  SDFF_X1 reg_out_reg_30_ ( .D(1'b0), .SI(n33), .SE(reg_in[30]), .CK(clk), .Q(
        reg_out[30]) );
  SDFF_X1 reg_out_reg_29_ ( .D(1'b0), .SI(n33), .SE(reg_in[29]), .CK(clk), .Q(
        reg_out[29]) );
  SDFF_X1 reg_out_reg_28_ ( .D(1'b0), .SI(n33), .SE(reg_in[28]), .CK(clk), .Q(
        reg_out[28]) );
  SDFF_X1 reg_out_reg_27_ ( .D(1'b0), .SI(n33), .SE(reg_in[27]), .CK(clk), .Q(
        reg_out[27]) );
  SDFF_X1 reg_out_reg_26_ ( .D(1'b0), .SI(n33), .SE(reg_in[26]), .CK(clk), .Q(
        reg_out[26]) );
  SDFF_X1 reg_out_reg_25_ ( .D(1'b0), .SI(n33), .SE(reg_in[25]), .CK(clk), .Q(
        reg_out[25]) );
  SDFF_X1 reg_out_reg_24_ ( .D(1'b0), .SI(n33), .SE(reg_in[24]), .CK(clk), .Q(
        reg_out[24]) );
  SDFF_X1 reg_out_reg_23_ ( .D(1'b0), .SI(n33), .SE(reg_in[23]), .CK(clk), .Q(
        reg_out[23]) );
  SDFF_X1 reg_out_reg_22_ ( .D(1'b0), .SI(n33), .SE(reg_in[22]), .CK(clk), .Q(
        reg_out[22]) );
  SDFF_X1 reg_out_reg_21_ ( .D(1'b0), .SI(n33), .SE(reg_in[21]), .CK(clk), .Q(
        reg_out[21]) );
  SDFF_X1 reg_out_reg_20_ ( .D(1'b0), .SI(n34), .SE(reg_in[20]), .CK(clk), .Q(
        reg_out[20]) );
  SDFF_X1 reg_out_reg_19_ ( .D(1'b0), .SI(n34), .SE(reg_in[19]), .CK(clk), .Q(
        reg_out[19]) );
  SDFF_X1 reg_out_reg_18_ ( .D(1'b0), .SI(n34), .SE(reg_in[18]), .CK(clk), .Q(
        reg_out[18]) );
  SDFF_X1 reg_out_reg_17_ ( .D(1'b0), .SI(n34), .SE(reg_in[17]), .CK(clk), .Q(
        reg_out[17]) );
  SDFF_X1 reg_out_reg_16_ ( .D(1'b0), .SI(n34), .SE(reg_in[16]), .CK(clk), .Q(
        reg_out[16]) );
  SDFF_X1 reg_out_reg_15_ ( .D(1'b0), .SI(n34), .SE(reg_in[15]), .CK(clk), .Q(
        reg_out[15]) );
  SDFF_X1 reg_out_reg_14_ ( .D(1'b0), .SI(n34), .SE(reg_in[14]), .CK(clk), .Q(
        reg_out[14]) );
  SDFF_X1 reg_out_reg_13_ ( .D(1'b0), .SI(n34), .SE(reg_in[13]), .CK(clk), .Q(
        reg_out[13]) );
  SDFF_X1 reg_out_reg_12_ ( .D(1'b0), .SI(n34), .SE(reg_in[12]), .CK(clk), .Q(
        reg_out[12]) );
  SDFF_X1 reg_out_reg_11_ ( .D(1'b0), .SI(n34), .SE(reg_in[11]), .CK(clk), .Q(
        reg_out[11]) );
  SDFF_X1 reg_out_reg_10_ ( .D(1'b0), .SI(n34), .SE(reg_in[10]), .CK(clk), .Q(
        reg_out[10]) );
  SDFF_X1 reg_out_reg_9_ ( .D(1'b0), .SI(n35), .SE(reg_in[9]), .CK(clk), .Q(
        reg_out[9]) );
  SDFF_X1 reg_out_reg_8_ ( .D(1'b0), .SI(n35), .SE(reg_in[8]), .CK(clk), .Q(
        reg_out[8]) );
  SDFF_X1 reg_out_reg_7_ ( .D(1'b0), .SI(n35), .SE(reg_in[7]), .CK(clk), .Q(
        reg_out[7]) );
  SDFF_X1 reg_out_reg_6_ ( .D(1'b0), .SI(n35), .SE(reg_in[6]), .CK(clk), .Q(
        reg_out[6]) );
  SDFF_X1 reg_out_reg_5_ ( .D(1'b0), .SI(n35), .SE(reg_in[5]), .CK(clk), .Q(
        reg_out[5]) );
  SDFF_X1 reg_out_reg_4_ ( .D(1'b0), .SI(n35), .SE(reg_in[4]), .CK(clk), .Q(
        reg_out[4]) );
  SDFF_X1 reg_out_reg_3_ ( .D(1'b0), .SI(n35), .SE(reg_in[3]), .CK(clk), .Q(
        reg_out[3]) );
  SDFF_X1 reg_out_reg_2_ ( .D(1'b0), .SI(n35), .SE(reg_in[2]), .CK(clk), .Q(
        reg_out[2]) );
  SDFF_X1 reg_out_reg_1_ ( .D(1'b0), .SI(n35), .SE(reg_in[1]), .CK(clk), .Q(
        reg_out[1]) );
  SDFF_X1 reg_out_reg_0_ ( .D(1'b0), .SI(n35), .SE(reg_in[0]), .CK(clk), .Q(
        reg_out[0]) );
  BUF_X1 U35 ( .A(n36), .Z(n34) );
  BUF_X1 U36 ( .A(n36), .Z(n33) );
  BUF_X1 U37 ( .A(n36), .Z(n35) );
  INV_X1 U38 ( .A(reset), .ZN(n36) );
endmodule


module simpleMultiplier_DW01_add_0 ( A, B, CI, SUM, CO );
  input [61:0] A;
  input [61:0] B;
  output [61:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180;
  assign SUM[29] = A[29];
  assign SUM[28] = A[28];
  assign SUM[27] = A[27];
  assign SUM[26] = A[26];
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .A(n110), .ZN(n25) );
  INV_X1 U3 ( .A(n107), .ZN(n23) );
  INV_X1 U4 ( .A(n144), .ZN(n27) );
  INV_X1 U5 ( .A(n131), .ZN(n21) );
  INV_X1 U6 ( .A(n111), .ZN(n14) );
  INV_X1 U7 ( .A(n88), .ZN(n12) );
  INV_X1 U8 ( .A(n80), .ZN(n10) );
  INV_X1 U9 ( .A(n72), .ZN(n8) );
  INV_X1 U10 ( .A(n64), .ZN(n6) );
  INV_X1 U11 ( .A(n56), .ZN(n4) );
  INV_X1 U12 ( .A(n48), .ZN(n2) );
  INV_X1 U13 ( .A(n145), .ZN(n29) );
  INV_X1 U14 ( .A(n172), .ZN(n35) );
  INV_X1 U15 ( .A(n142), .ZN(n26) );
  INV_X1 U16 ( .A(n50), .ZN(n3) );
  INV_X1 U17 ( .A(n42), .ZN(n1) );
  INV_X1 U18 ( .A(n149), .ZN(n31) );
  INV_X1 U19 ( .A(n127), .ZN(n20) );
  INV_X1 U20 ( .A(n122), .ZN(n18) );
  INV_X1 U21 ( .A(n102), .ZN(n17) );
  INV_X1 U22 ( .A(n97), .ZN(n15) );
  INV_X1 U23 ( .A(n90), .ZN(n13) );
  INV_X1 U24 ( .A(n82), .ZN(n11) );
  INV_X1 U25 ( .A(n74), .ZN(n9) );
  INV_X1 U26 ( .A(n66), .ZN(n7) );
  INV_X1 U27 ( .A(n58), .ZN(n5) );
  INV_X1 U28 ( .A(n158), .ZN(n34) );
  INV_X1 U29 ( .A(n165), .ZN(n36) );
  INV_X1 U30 ( .A(n106), .ZN(n24) );
  INV_X1 U31 ( .A(n130), .ZN(n19) );
  INV_X1 U32 ( .A(n148), .ZN(n28) );
  INV_X1 U33 ( .A(n170), .ZN(n33) );
  INV_X1 U34 ( .A(n160), .ZN(n32) );
  INV_X1 U35 ( .A(n117), .ZN(n16) );
  INV_X1 U36 ( .A(n147), .ZN(n30) );
  INV_X1 U37 ( .A(n128), .ZN(n22) );
  INV_X1 U38 ( .A(n176), .ZN(n38) );
  INV_X1 U39 ( .A(n175), .ZN(n37) );
  INV_X1 U40 ( .A(n180), .ZN(SUM[30]) );
  XOR2_X1 U41 ( .A(n40), .B(n41), .Z(SUM[61]) );
  XOR2_X1 U42 ( .A(B[61]), .B(A[61]), .Z(n41) );
  OAI21_X1 U43 ( .B1(n42), .B2(n43), .A(n44), .ZN(n40) );
  XOR2_X1 U44 ( .A(n45), .B(n43), .Z(SUM[60]) );
  AOI21_X1 U45 ( .B1(n2), .B2(n46), .A(n47), .ZN(n43) );
  NAND2_X1 U46 ( .A1(n1), .A2(n44), .ZN(n45) );
  NAND2_X1 U47 ( .A1(B[60]), .A2(A[60]), .ZN(n44) );
  NOR2_X1 U48 ( .A1(B[60]), .A2(A[60]), .ZN(n42) );
  XOR2_X1 U49 ( .A(n46), .B(n49), .Z(SUM[59]) );
  NOR2_X1 U50 ( .A1(n47), .A2(n48), .ZN(n49) );
  NOR2_X1 U51 ( .A1(B[59]), .A2(A[59]), .ZN(n48) );
  AND2_X1 U52 ( .A1(B[59]), .A2(A[59]), .ZN(n47) );
  OAI21_X1 U53 ( .B1(n50), .B2(n51), .A(n52), .ZN(n46) );
  XOR2_X1 U54 ( .A(n53), .B(n51), .Z(SUM[58]) );
  AOI21_X1 U55 ( .B1(n4), .B2(n54), .A(n55), .ZN(n51) );
  NAND2_X1 U56 ( .A1(n3), .A2(n52), .ZN(n53) );
  NAND2_X1 U57 ( .A1(B[58]), .A2(A[58]), .ZN(n52) );
  NOR2_X1 U58 ( .A1(B[58]), .A2(A[58]), .ZN(n50) );
  XOR2_X1 U59 ( .A(n54), .B(n57), .Z(SUM[57]) );
  NOR2_X1 U60 ( .A1(n55), .A2(n56), .ZN(n57) );
  NOR2_X1 U61 ( .A1(B[57]), .A2(A[57]), .ZN(n56) );
  AND2_X1 U62 ( .A1(B[57]), .A2(A[57]), .ZN(n55) );
  OAI21_X1 U63 ( .B1(n58), .B2(n59), .A(n60), .ZN(n54) );
  XOR2_X1 U64 ( .A(n61), .B(n59), .Z(SUM[56]) );
  AOI21_X1 U65 ( .B1(n6), .B2(n62), .A(n63), .ZN(n59) );
  NAND2_X1 U66 ( .A1(n5), .A2(n60), .ZN(n61) );
  NAND2_X1 U67 ( .A1(B[56]), .A2(A[56]), .ZN(n60) );
  NOR2_X1 U68 ( .A1(B[56]), .A2(A[56]), .ZN(n58) );
  XOR2_X1 U69 ( .A(n62), .B(n65), .Z(SUM[55]) );
  NOR2_X1 U70 ( .A1(n63), .A2(n64), .ZN(n65) );
  NOR2_X1 U71 ( .A1(B[55]), .A2(A[55]), .ZN(n64) );
  AND2_X1 U72 ( .A1(B[55]), .A2(A[55]), .ZN(n63) );
  OAI21_X1 U73 ( .B1(n66), .B2(n67), .A(n68), .ZN(n62) );
  XOR2_X1 U74 ( .A(n69), .B(n67), .Z(SUM[54]) );
  AOI21_X1 U75 ( .B1(n8), .B2(n70), .A(n71), .ZN(n67) );
  NAND2_X1 U76 ( .A1(n7), .A2(n68), .ZN(n69) );
  NAND2_X1 U77 ( .A1(B[54]), .A2(A[54]), .ZN(n68) );
  NOR2_X1 U78 ( .A1(B[54]), .A2(A[54]), .ZN(n66) );
  XOR2_X1 U79 ( .A(n70), .B(n73), .Z(SUM[53]) );
  NOR2_X1 U80 ( .A1(n71), .A2(n72), .ZN(n73) );
  NOR2_X1 U81 ( .A1(B[53]), .A2(A[53]), .ZN(n72) );
  AND2_X1 U82 ( .A1(B[53]), .A2(A[53]), .ZN(n71) );
  OAI21_X1 U83 ( .B1(n74), .B2(n75), .A(n76), .ZN(n70) );
  XOR2_X1 U84 ( .A(n77), .B(n75), .Z(SUM[52]) );
  AOI21_X1 U85 ( .B1(n10), .B2(n78), .A(n79), .ZN(n75) );
  NAND2_X1 U86 ( .A1(n9), .A2(n76), .ZN(n77) );
  NAND2_X1 U87 ( .A1(B[52]), .A2(A[52]), .ZN(n76) );
  NOR2_X1 U88 ( .A1(B[52]), .A2(A[52]), .ZN(n74) );
  XOR2_X1 U89 ( .A(n78), .B(n81), .Z(SUM[51]) );
  NOR2_X1 U90 ( .A1(n79), .A2(n80), .ZN(n81) );
  NOR2_X1 U91 ( .A1(B[51]), .A2(A[51]), .ZN(n80) );
  AND2_X1 U92 ( .A1(B[51]), .A2(A[51]), .ZN(n79) );
  OAI21_X1 U93 ( .B1(n82), .B2(n83), .A(n84), .ZN(n78) );
  XOR2_X1 U94 ( .A(n85), .B(n83), .Z(SUM[50]) );
  AOI21_X1 U95 ( .B1(n12), .B2(n86), .A(n87), .ZN(n83) );
  NAND2_X1 U96 ( .A1(n11), .A2(n84), .ZN(n85) );
  NAND2_X1 U97 ( .A1(B[50]), .A2(A[50]), .ZN(n84) );
  NOR2_X1 U98 ( .A1(B[50]), .A2(A[50]), .ZN(n82) );
  XOR2_X1 U99 ( .A(n86), .B(n89), .Z(SUM[49]) );
  NOR2_X1 U100 ( .A1(n87), .A2(n88), .ZN(n89) );
  NOR2_X1 U101 ( .A1(B[49]), .A2(A[49]), .ZN(n88) );
  AND2_X1 U102 ( .A1(B[49]), .A2(A[49]), .ZN(n87) );
  OAI21_X1 U103 ( .B1(n90), .B2(n91), .A(n92), .ZN(n86) );
  XOR2_X1 U104 ( .A(n93), .B(n91), .Z(SUM[48]) );
  AOI21_X1 U105 ( .B1(n14), .B2(n94), .A(n95), .ZN(n91) );
  OAI21_X1 U106 ( .B1(n96), .B2(n97), .A(n98), .ZN(n94) );
  AOI21_X1 U107 ( .B1(n16), .B2(n99), .A(n100), .ZN(n96) );
  OAI21_X1 U108 ( .B1(n101), .B2(n102), .A(n103), .ZN(n99) );
  AOI21_X1 U109 ( .B1(n24), .B2(n104), .A(n105), .ZN(n101) );
  AOI221_X1 U110 ( .B1(n107), .B2(n108), .C1(n109), .C2(n107), .A(n110), .ZN(
        n106) );
  NAND2_X1 U111 ( .A1(n13), .A2(n92), .ZN(n93) );
  NAND2_X1 U112 ( .A1(B[48]), .A2(A[48]), .ZN(n92) );
  NOR2_X1 U113 ( .A1(B[48]), .A2(A[48]), .ZN(n90) );
  XOR2_X1 U114 ( .A(n112), .B(n113), .Z(SUM[47]) );
  NOR2_X1 U115 ( .A1(n95), .A2(n111), .ZN(n113) );
  NOR2_X1 U116 ( .A1(B[47]), .A2(A[47]), .ZN(n111) );
  AND2_X1 U117 ( .A1(B[47]), .A2(A[47]), .ZN(n95) );
  OAI21_X1 U118 ( .B1(n97), .B2(n114), .A(n98), .ZN(n112) );
  XOR2_X1 U119 ( .A(n115), .B(n114), .Z(SUM[46]) );
  AOI21_X1 U120 ( .B1(n16), .B2(n116), .A(n100), .ZN(n114) );
  NAND2_X1 U121 ( .A1(n15), .A2(n98), .ZN(n115) );
  NAND2_X1 U122 ( .A1(B[46]), .A2(A[46]), .ZN(n98) );
  NOR2_X1 U123 ( .A1(B[46]), .A2(A[46]), .ZN(n97) );
  XOR2_X1 U124 ( .A(n116), .B(n118), .Z(SUM[45]) );
  NOR2_X1 U125 ( .A1(n100), .A2(n117), .ZN(n118) );
  NOR2_X1 U126 ( .A1(B[45]), .A2(A[45]), .ZN(n117) );
  AND2_X1 U127 ( .A1(B[45]), .A2(A[45]), .ZN(n100) );
  OAI21_X1 U128 ( .B1(n102), .B2(n119), .A(n103), .ZN(n116) );
  XOR2_X1 U129 ( .A(n120), .B(n119), .Z(SUM[44]) );
  AOI21_X1 U130 ( .B1(n121), .B2(n104), .A(n105), .ZN(n119) );
  OAI21_X1 U131 ( .B1(n122), .B2(n123), .A(n124), .ZN(n105) );
  AOI21_X1 U132 ( .B1(n125), .B2(n19), .A(n126), .ZN(n123) );
  OAI21_X1 U133 ( .B1(n127), .B2(n128), .A(n129), .ZN(n125) );
  NOR4_X1 U134 ( .A1(n122), .A2(n130), .A3(n127), .A4(n131), .ZN(n104) );
  NAND2_X1 U135 ( .A1(n17), .A2(n103), .ZN(n120) );
  NAND2_X1 U136 ( .A1(B[44]), .A2(A[44]), .ZN(n103) );
  NOR2_X1 U137 ( .A1(B[44]), .A2(A[44]), .ZN(n102) );
  XOR2_X1 U138 ( .A(n132), .B(n133), .Z(SUM[43]) );
  AOI21_X1 U139 ( .B1(n134), .B2(n19), .A(n126), .ZN(n133) );
  NAND2_X1 U140 ( .A1(n18), .A2(n124), .ZN(n132) );
  NAND2_X1 U141 ( .A1(B[43]), .A2(A[43]), .ZN(n124) );
  NOR2_X1 U142 ( .A1(B[43]), .A2(A[43]), .ZN(n122) );
  XOR2_X1 U143 ( .A(n134), .B(n135), .Z(SUM[42]) );
  NOR2_X1 U144 ( .A1(n126), .A2(n130), .ZN(n135) );
  NOR2_X1 U145 ( .A1(B[42]), .A2(A[42]), .ZN(n130) );
  AND2_X1 U146 ( .A1(B[42]), .A2(A[42]), .ZN(n126) );
  OAI21_X1 U147 ( .B1(n127), .B2(n136), .A(n129), .ZN(n134) );
  XOR2_X1 U148 ( .A(n137), .B(n136), .Z(SUM[41]) );
  AOI21_X1 U149 ( .B1(n21), .B2(n121), .A(n22), .ZN(n136) );
  NAND2_X1 U150 ( .A1(n20), .A2(n129), .ZN(n137) );
  NAND2_X1 U151 ( .A1(B[41]), .A2(A[41]), .ZN(n129) );
  NOR2_X1 U152 ( .A1(B[41]), .A2(A[41]), .ZN(n127) );
  XOR2_X1 U153 ( .A(n121), .B(n138), .Z(SUM[40]) );
  NOR2_X1 U154 ( .A1(n22), .A2(n131), .ZN(n138) );
  NOR2_X1 U155 ( .A1(B[40]), .A2(A[40]), .ZN(n131) );
  NAND2_X1 U156 ( .A1(B[40]), .A2(A[40]), .ZN(n128) );
  OAI21_X1 U157 ( .B1(n139), .B2(n23), .A(n25), .ZN(n121) );
  OAI21_X1 U158 ( .B1(n140), .B2(n141), .A(n142), .ZN(n110) );
  AOI21_X1 U159 ( .B1(n143), .B2(n28), .A(n27), .ZN(n141) );
  OAI21_X1 U160 ( .B1(n145), .B2(n146), .A(n147), .ZN(n143) );
  NOR4_X1 U161 ( .A1(n140), .A2(n148), .A3(n145), .A4(n149), .ZN(n107) );
  XOR2_X1 U162 ( .A(n150), .B(n151), .Z(SUM[39]) );
  NOR2_X1 U163 ( .A1(n26), .A2(n140), .ZN(n151) );
  NOR2_X1 U164 ( .A1(B[39]), .A2(A[39]), .ZN(n140) );
  NAND2_X1 U165 ( .A1(B[39]), .A2(A[39]), .ZN(n142) );
  OAI21_X1 U166 ( .B1(n148), .B2(n152), .A(n144), .ZN(n150) );
  XOR2_X1 U167 ( .A(n153), .B(n152), .Z(SUM[38]) );
  AOI21_X1 U168 ( .B1(n29), .B2(n154), .A(n30), .ZN(n152) );
  NAND2_X1 U169 ( .A1(n28), .A2(n144), .ZN(n153) );
  NAND2_X1 U170 ( .A1(B[38]), .A2(A[38]), .ZN(n144) );
  NOR2_X1 U171 ( .A1(B[38]), .A2(A[38]), .ZN(n148) );
  XOR2_X1 U172 ( .A(n154), .B(n155), .Z(SUM[37]) );
  NOR2_X1 U173 ( .A1(n30), .A2(n145), .ZN(n155) );
  NOR2_X1 U174 ( .A1(B[37]), .A2(A[37]), .ZN(n145) );
  NAND2_X1 U175 ( .A1(B[37]), .A2(A[37]), .ZN(n147) );
  OAI21_X1 U176 ( .B1(n149), .B2(n139), .A(n146), .ZN(n154) );
  XOR2_X1 U177 ( .A(n156), .B(n139), .Z(SUM[36]) );
  NOR2_X1 U178 ( .A1(n108), .A2(n109), .ZN(n139) );
  NOR4_X1 U179 ( .A1(n37), .A2(n157), .A3(n158), .A4(n159), .ZN(n109) );
  NAND2_X1 U180 ( .A1(n33), .A2(n32), .ZN(n159) );
  OAI21_X1 U181 ( .B1(n160), .B2(n161), .A(n162), .ZN(n108) );
  AOI21_X1 U182 ( .B1(n163), .B2(n33), .A(n164), .ZN(n161) );
  OAI21_X1 U183 ( .B1(n158), .B2(n165), .A(n166), .ZN(n163) );
  NAND2_X1 U184 ( .A1(n31), .A2(n146), .ZN(n156) );
  NAND2_X1 U185 ( .A1(B[36]), .A2(A[36]), .ZN(n146) );
  NOR2_X1 U186 ( .A1(B[36]), .A2(A[36]), .ZN(n149) );
  XOR2_X1 U187 ( .A(n167), .B(n168), .Z(SUM[35]) );
  AOI21_X1 U188 ( .B1(n169), .B2(n33), .A(n164), .ZN(n168) );
  NAND2_X1 U189 ( .A1(n32), .A2(n162), .ZN(n167) );
  NAND2_X1 U190 ( .A1(B[35]), .A2(A[35]), .ZN(n162) );
  NOR2_X1 U191 ( .A1(B[35]), .A2(A[35]), .ZN(n160) );
  XOR2_X1 U192 ( .A(n169), .B(n171), .Z(SUM[34]) );
  NOR2_X1 U193 ( .A1(n164), .A2(n170), .ZN(n171) );
  NOR2_X1 U194 ( .A1(B[34]), .A2(A[34]), .ZN(n170) );
  AND2_X1 U195 ( .A1(B[34]), .A2(A[34]), .ZN(n164) );
  OAI21_X1 U196 ( .B1(n158), .B2(n35), .A(n166), .ZN(n169) );
  XNOR2_X1 U197 ( .A(n173), .B(n172), .ZN(SUM[33]) );
  OAI21_X1 U198 ( .B1(n157), .B2(n37), .A(n165), .ZN(n172) );
  NAND2_X1 U199 ( .A1(n34), .A2(n166), .ZN(n173) );
  NAND2_X1 U200 ( .A1(B[33]), .A2(A[33]), .ZN(n166) );
  NOR2_X1 U201 ( .A1(B[33]), .A2(A[33]), .ZN(n158) );
  XNOR2_X1 U202 ( .A(n37), .B(n174), .ZN(SUM[32]) );
  NOR2_X1 U203 ( .A1(n36), .A2(n157), .ZN(n174) );
  NOR2_X1 U204 ( .A1(B[32]), .A2(A[32]), .ZN(n157) );
  NAND2_X1 U205 ( .A1(B[32]), .A2(A[32]), .ZN(n165) );
  OAI21_X1 U206 ( .B1(n176), .B2(n177), .A(n178), .ZN(n175) );
  XOR2_X1 U207 ( .A(n177), .B(n179), .Z(SUM[31]) );
  NAND2_X1 U208 ( .A1(n38), .A2(n178), .ZN(n179) );
  NAND2_X1 U209 ( .A1(B[31]), .A2(A[31]), .ZN(n178) );
  NOR2_X1 U210 ( .A1(B[31]), .A2(A[31]), .ZN(n176) );
  OAI21_X1 U211 ( .B1(B[30]), .B2(A[30]), .A(n177), .ZN(n180) );
  NAND2_X1 U212 ( .A1(B[30]), .A2(A[30]), .ZN(n177) );
endmodule


module simpleMultiplier_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   ab_31__31_, ab_31__30_, ab_31__29_, ab_31__28_, ab_31__27_,
         ab_31__26_, ab_31__25_, ab_31__24_, ab_31__23_, ab_31__22_,
         ab_31__21_, ab_31__20_, ab_31__19_, ab_31__18_, ab_31__17_,
         ab_31__16_, ab_31__15_, ab_31__14_, ab_31__13_, ab_31__12_,
         ab_31__11_, ab_31__10_, ab_31__9_, ab_31__8_, ab_31__7_, ab_31__6_,
         ab_31__5_, ab_31__4_, ab_31__3_, ab_31__2_, ab_31__1_, ab_31__0_,
         ab_30__31_, ab_30__30_, ab_30__29_, ab_30__28_, ab_30__27_,
         ab_30__26_, ab_30__25_, ab_30__24_, ab_30__23_, ab_30__22_,
         ab_30__21_, ab_30__20_, ab_30__19_, ab_30__18_, ab_30__17_,
         ab_30__16_, ab_30__15_, ab_30__14_, ab_30__13_, ab_30__12_,
         ab_30__11_, ab_30__10_, ab_30__9_, ab_30__8_, ab_30__7_, ab_30__6_,
         ab_30__5_, ab_30__4_, ab_30__3_, ab_30__2_, ab_30__1_, ab_30__0_,
         ab_29__31_, ab_29__30_, ab_29__29_, ab_29__28_, ab_29__27_,
         ab_29__26_, ab_29__25_, ab_29__24_, ab_29__23_, ab_29__22_,
         ab_29__21_, ab_29__20_, ab_29__19_, ab_29__18_, ab_29__17_,
         ab_29__16_, ab_29__15_, ab_29__14_, ab_29__13_, ab_29__12_,
         ab_29__11_, ab_29__10_, ab_29__9_, ab_29__8_, ab_29__7_, ab_29__6_,
         ab_29__5_, ab_29__4_, ab_29__3_, ab_29__2_, ab_29__1_, ab_29__0_,
         ab_28__31_, ab_28__30_, ab_28__29_, ab_28__28_, ab_28__27_,
         ab_28__26_, ab_28__25_, ab_28__24_, ab_28__23_, ab_28__22_,
         ab_28__21_, ab_28__20_, ab_28__19_, ab_28__18_, ab_28__17_,
         ab_28__16_, ab_28__15_, ab_28__14_, ab_28__13_, ab_28__12_,
         ab_28__11_, ab_28__10_, ab_28__9_, ab_28__8_, ab_28__7_, ab_28__6_,
         ab_28__5_, ab_28__4_, ab_28__3_, ab_28__2_, ab_28__1_, ab_28__0_,
         ab_27__31_, ab_27__30_, ab_27__29_, ab_27__28_, ab_27__27_,
         ab_27__26_, ab_27__25_, ab_27__24_, ab_27__23_, ab_27__22_,
         ab_27__21_, ab_27__20_, ab_27__19_, ab_27__18_, ab_27__17_,
         ab_27__16_, ab_27__15_, ab_27__14_, ab_27__13_, ab_27__12_,
         ab_27__11_, ab_27__10_, ab_27__9_, ab_27__8_, ab_27__7_, ab_27__6_,
         ab_27__5_, ab_27__4_, ab_27__3_, ab_27__2_, ab_27__1_, ab_27__0_,
         ab_26__31_, ab_26__30_, ab_26__29_, ab_26__28_, ab_26__27_,
         ab_26__26_, ab_26__25_, ab_26__24_, ab_26__23_, ab_26__22_,
         ab_26__21_, ab_26__20_, ab_26__19_, ab_26__18_, ab_26__17_,
         ab_26__16_, ab_26__15_, ab_26__14_, ab_26__13_, ab_26__12_,
         ab_26__11_, ab_26__10_, ab_26__9_, ab_26__8_, ab_26__7_, ab_26__6_,
         ab_26__5_, ab_26__4_, ab_26__3_, ab_26__2_, ab_26__1_, ab_26__0_,
         ab_25__31_, ab_25__30_, ab_25__29_, ab_25__28_, ab_25__27_,
         ab_25__26_, ab_25__25_, ab_25__24_, ab_25__23_, ab_25__22_,
         ab_25__21_, ab_25__20_, ab_25__19_, ab_25__18_, ab_25__17_,
         ab_25__16_, ab_25__15_, ab_25__14_, ab_25__13_, ab_25__12_,
         ab_25__11_, ab_25__10_, ab_25__9_, ab_25__8_, ab_25__7_, ab_25__6_,
         ab_25__5_, ab_25__4_, ab_25__3_, ab_25__2_, ab_25__1_, ab_25__0_,
         ab_24__31_, ab_24__30_, ab_24__29_, ab_24__28_, ab_24__27_,
         ab_24__26_, ab_24__25_, ab_24__24_, ab_24__23_, ab_24__22_,
         ab_24__21_, ab_24__20_, ab_24__19_, ab_24__18_, ab_24__17_,
         ab_24__16_, ab_24__15_, ab_24__14_, ab_24__13_, ab_24__12_,
         ab_24__11_, ab_24__10_, ab_24__9_, ab_24__8_, ab_24__7_, ab_24__6_,
         ab_24__5_, ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_,
         ab_23__31_, ab_23__30_, ab_23__29_, ab_23__28_, ab_23__27_,
         ab_23__26_, ab_23__25_, ab_23__24_, ab_23__23_, ab_23__22_,
         ab_23__21_, ab_23__20_, ab_23__19_, ab_23__18_, ab_23__17_,
         ab_23__16_, ab_23__15_, ab_23__14_, ab_23__13_, ab_23__12_,
         ab_23__11_, ab_23__10_, ab_23__9_, ab_23__8_, ab_23__7_, ab_23__6_,
         ab_23__5_, ab_23__4_, ab_23__3_, ab_23__2_, ab_23__1_, ab_23__0_,
         ab_22__31_, ab_22__30_, ab_22__29_, ab_22__28_, ab_22__27_,
         ab_22__26_, ab_22__25_, ab_22__24_, ab_22__23_, ab_22__22_,
         ab_22__21_, ab_22__20_, ab_22__19_, ab_22__18_, ab_22__17_,
         ab_22__16_, ab_22__15_, ab_22__14_, ab_22__13_, ab_22__12_,
         ab_22__11_, ab_22__10_, ab_22__9_, ab_22__8_, ab_22__7_, ab_22__6_,
         ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_, ab_22__0_,
         ab_21__31_, ab_21__30_, ab_21__29_, ab_21__28_, ab_21__27_,
         ab_21__26_, ab_21__25_, ab_21__24_, ab_21__23_, ab_21__22_,
         ab_21__21_, ab_21__20_, ab_21__19_, ab_21__18_, ab_21__17_,
         ab_21__16_, ab_21__15_, ab_21__14_, ab_21__13_, ab_21__12_,
         ab_21__11_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_,
         ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_,
         ab_20__31_, ab_20__30_, ab_20__29_, ab_20__28_, ab_20__27_,
         ab_20__26_, ab_20__25_, ab_20__24_, ab_20__23_, ab_20__22_,
         ab_20__21_, ab_20__20_, ab_20__19_, ab_20__18_, ab_20__17_,
         ab_20__16_, ab_20__15_, ab_20__14_, ab_20__13_, ab_20__12_,
         ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_,
         ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_,
         ab_19__31_, ab_19__30_, ab_19__29_, ab_19__28_, ab_19__27_,
         ab_19__26_, ab_19__25_, ab_19__24_, ab_19__23_, ab_19__22_,
         ab_19__21_, ab_19__20_, ab_19__19_, ab_19__18_, ab_19__17_,
         ab_19__16_, ab_19__15_, ab_19__14_, ab_19__13_, ab_19__12_,
         ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_, ab_19__6_,
         ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_, ab_19__0_,
         ab_18__31_, ab_18__30_, ab_18__29_, ab_18__28_, ab_18__27_,
         ab_18__26_, ab_18__25_, ab_18__24_, ab_18__23_, ab_18__22_,
         ab_18__21_, ab_18__20_, ab_18__19_, ab_18__18_, ab_18__17_,
         ab_18__16_, ab_18__15_, ab_18__14_, ab_18__13_, ab_18__12_,
         ab_18__11_, ab_18__10_, ab_18__9_, ab_18__8_, ab_18__7_, ab_18__6_,
         ab_18__5_, ab_18__4_, ab_18__3_, ab_18__2_, ab_18__1_, ab_18__0_,
         ab_17__31_, ab_17__30_, ab_17__29_, ab_17__28_, ab_17__27_,
         ab_17__26_, ab_17__25_, ab_17__24_, ab_17__23_, ab_17__22_,
         ab_17__21_, ab_17__20_, ab_17__19_, ab_17__18_, ab_17__17_,
         ab_17__16_, ab_17__15_, ab_17__14_, ab_17__13_, ab_17__12_,
         ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_,
         ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_,
         ab_16__31_, ab_16__30_, ab_16__29_, ab_16__28_, ab_16__27_,
         ab_16__26_, ab_16__25_, ab_16__24_, ab_16__23_, ab_16__22_,
         ab_16__21_, ab_16__20_, ab_16__19_, ab_16__18_, ab_16__17_,
         ab_16__16_, ab_16__15_, ab_16__14_, ab_16__13_, ab_16__12_,
         ab_16__11_, ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_, ab_16__6_,
         ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_, ab_16__0_,
         ab_15__31_, ab_15__30_, ab_15__29_, ab_15__28_, ab_15__27_,
         ab_15__26_, ab_15__25_, ab_15__24_, ab_15__23_, ab_15__22_,
         ab_15__21_, ab_15__20_, ab_15__19_, ab_15__18_, ab_15__17_,
         ab_15__16_, ab_15__15_, ab_15__14_, ab_15__13_, ab_15__12_,
         ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_, ab_15__6_,
         ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_,
         ab_14__31_, ab_14__30_, ab_14__29_, ab_14__28_, ab_14__27_,
         ab_14__26_, ab_14__25_, ab_14__24_, ab_14__23_, ab_14__22_,
         ab_14__21_, ab_14__20_, ab_14__19_, ab_14__18_, ab_14__17_,
         ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__31_, ab_13__30_, ab_13__29_, ab_13__28_, ab_13__27_,
         ab_13__26_, ab_13__25_, ab_13__24_, ab_13__23_, ab_13__22_,
         ab_13__21_, ab_13__20_, ab_13__19_, ab_13__18_, ab_13__17_,
         ab_13__16_, ab_13__15_, ab_13__14_, ab_13__13_, ab_13__12_,
         ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_, ab_13__6_,
         ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_, ab_13__0_,
         ab_12__31_, ab_12__30_, ab_12__29_, ab_12__28_, ab_12__27_,
         ab_12__26_, ab_12__25_, ab_12__24_, ab_12__23_, ab_12__22_,
         ab_12__21_, ab_12__20_, ab_12__19_, ab_12__18_, ab_12__17_,
         ab_12__16_, ab_12__15_, ab_12__14_, ab_12__13_, ab_12__12_,
         ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_, ab_12__6_,
         ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_,
         ab_11__31_, ab_11__30_, ab_11__29_, ab_11__28_, ab_11__27_,
         ab_11__26_, ab_11__25_, ab_11__24_, ab_11__23_, ab_11__22_,
         ab_11__21_, ab_11__20_, ab_11__19_, ab_11__18_, ab_11__17_,
         ab_11__16_, ab_11__15_, ab_11__14_, ab_11__13_, ab_11__12_,
         ab_11__11_, ab_11__10_, ab_11__9_, ab_11__8_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__31_, ab_10__30_, ab_10__29_, ab_10__28_, ab_10__27_,
         ab_10__26_, ab_10__25_, ab_10__24_, ab_10__23_, ab_10__22_,
         ab_10__21_, ab_10__20_, ab_10__19_, ab_10__18_, ab_10__17_,
         ab_10__16_, ab_10__15_, ab_10__14_, ab_10__13_, ab_10__12_,
         ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_, ab_10__7_, ab_10__6_,
         ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_, ab_10__1_, ab_10__0_,
         ab_9__31_, ab_9__30_, ab_9__29_, ab_9__28_, ab_9__27_, ab_9__26_,
         ab_9__25_, ab_9__24_, ab_9__23_, ab_9__22_, ab_9__21_, ab_9__20_,
         ab_9__19_, ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_,
         ab_9__13_, ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_,
         ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_,
         ab_9__0_, ab_8__31_, ab_8__30_, ab_8__29_, ab_8__28_, ab_8__27_,
         ab_8__26_, ab_8__25_, ab_8__24_, ab_8__23_, ab_8__22_, ab_8__21_,
         ab_8__20_, ab_8__19_, ab_8__18_, ab_8__17_, ab_8__16_, ab_8__15_,
         ab_8__14_, ab_8__13_, ab_8__12_, ab_8__11_, ab_8__10_, ab_8__9_,
         ab_8__8_, ab_8__7_, ab_8__6_, ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_,
         ab_8__1_, ab_8__0_, ab_7__31_, ab_7__30_, ab_7__29_, ab_7__28_,
         ab_7__27_, ab_7__26_, ab_7__25_, ab_7__24_, ab_7__23_, ab_7__22_,
         ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_, ab_7__17_, ab_7__16_,
         ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_, ab_7__11_, ab_7__10_,
         ab_7__9_, ab_7__8_, ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_,
         ab_7__2_, ab_7__1_, ab_7__0_, ab_6__31_, ab_6__30_, ab_6__29_,
         ab_6__28_, ab_6__27_, ab_6__26_, ab_6__25_, ab_6__24_, ab_6__23_,
         ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_, ab_6__18_, ab_6__17_,
         ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_, ab_6__12_, ab_6__11_,
         ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_,
         ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_, ab_5__31_, ab_5__30_,
         ab_5__29_, ab_5__28_, ab_5__27_, ab_5__26_, ab_5__25_, ab_5__24_,
         ab_5__23_, ab_5__22_, ab_5__21_, ab_5__20_, ab_5__19_, ab_5__18_,
         ab_5__17_, ab_5__16_, ab_5__15_, ab_5__14_, ab_5__13_, ab_5__12_,
         ab_5__11_, ab_5__10_, ab_5__9_, ab_5__8_, ab_5__7_, ab_5__6_,
         ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_, ab_5__0_, ab_4__31_,
         ab_4__30_, ab_4__29_, ab_4__28_, ab_4__27_, ab_4__26_, ab_4__25_,
         ab_4__24_, ab_4__23_, ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_,
         ab_4__18_, ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_,
         ab_4__12_, ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_, ab_4__7_,
         ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_,
         ab_3__31_, ab_3__30_, ab_3__29_, ab_3__28_, ab_3__27_, ab_3__26_,
         ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_, ab_3__21_, ab_3__20_,
         ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_, ab_3__15_, ab_3__14_,
         ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_, ab_3__9_, ab_3__8_,
         ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_,
         ab_3__0_, ab_2__31_, ab_2__30_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_,
         ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_,
         ab_2__1_, ab_2__0_, ab_1__31_, ab_1__30_, ab_1__29_, ab_1__28_,
         ab_1__27_, ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_,
         ab_1__21_, ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_,
         ab_1__15_, ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_,
         ab_1__9_, ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_,
         ab_1__2_, ab_1__1_, ab_1__0_, ab_0__31_, ab_0__30_, ab_0__29_,
         ab_0__28_, ab_0__27_, ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_,
         ab_0__22_, ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_,
         ab_0__16_, ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_,
         ab_0__10_, ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, ab_0__1_, CARRYB_15__30_, CARRYB_15__29_,
         CARRYB_15__28_, CARRYB_15__27_, CARRYB_15__26_, CARRYB_15__25_,
         CARRYB_15__24_, CARRYB_15__23_, CARRYB_15__22_, CARRYB_15__21_,
         CARRYB_15__20_, CARRYB_15__19_, CARRYB_15__18_, CARRYB_15__17_,
         CARRYB_15__16_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__30_, CARRYB_14__29_, CARRYB_14__28_,
         CARRYB_14__27_, CARRYB_14__26_, CARRYB_14__25_, CARRYB_14__24_,
         CARRYB_14__23_, CARRYB_14__22_, CARRYB_14__21_, CARRYB_14__20_,
         CARRYB_14__19_, CARRYB_14__18_, CARRYB_14__17_, CARRYB_14__16_,
         CARRYB_14__15_, CARRYB_14__14_, CARRYB_14__13_, CARRYB_14__12_,
         CARRYB_14__11_, CARRYB_14__10_, CARRYB_14__9_, CARRYB_14__8_,
         CARRYB_14__7_, CARRYB_14__6_, CARRYB_14__5_, CARRYB_14__4_,
         CARRYB_14__3_, CARRYB_14__2_, CARRYB_14__1_, CARRYB_14__0_,
         CARRYB_13__30_, CARRYB_13__29_, CARRYB_13__28_, CARRYB_13__27_,
         CARRYB_13__26_, CARRYB_13__25_, CARRYB_13__24_, CARRYB_13__23_,
         CARRYB_13__22_, CARRYB_13__21_, CARRYB_13__20_, CARRYB_13__19_,
         CARRYB_13__18_, CARRYB_13__17_, CARRYB_13__16_, CARRYB_13__15_,
         CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_, CARRYB_13__11_,
         CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_, CARRYB_13__7_,
         CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_, CARRYB_13__3_,
         CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_, CARRYB_12__30_,
         CARRYB_12__29_, CARRYB_12__28_, CARRYB_12__27_, CARRYB_12__26_,
         CARRYB_12__25_, CARRYB_12__24_, CARRYB_12__23_, CARRYB_12__22_,
         CARRYB_12__21_, CARRYB_12__20_, CARRYB_12__19_, CARRYB_12__18_,
         CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_, CARRYB_12__14_,
         CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_, CARRYB_12__10_,
         CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_, CARRYB_12__6_,
         CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_, CARRYB_12__2_,
         CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__30_, CARRYB_11__29_,
         CARRYB_11__28_, CARRYB_11__27_, CARRYB_11__26_, CARRYB_11__25_,
         CARRYB_11__24_, CARRYB_11__23_, CARRYB_11__22_, CARRYB_11__21_,
         CARRYB_11__20_, CARRYB_11__19_, CARRYB_11__18_, CARRYB_11__17_,
         CARRYB_11__16_, CARRYB_11__15_, CARRYB_11__14_, CARRYB_11__13_,
         CARRYB_11__12_, CARRYB_11__11_, CARRYB_11__10_, CARRYB_11__9_,
         CARRYB_11__8_, CARRYB_11__7_, CARRYB_11__6_, CARRYB_11__5_,
         CARRYB_11__4_, CARRYB_11__3_, CARRYB_11__2_, CARRYB_11__1_,
         CARRYB_11__0_, CARRYB_10__30_, CARRYB_10__29_, CARRYB_10__28_,
         CARRYB_10__27_, CARRYB_10__26_, CARRYB_10__25_, CARRYB_10__24_,
         CARRYB_10__23_, CARRYB_10__22_, CARRYB_10__21_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__30_, CARRYB_9__29_, CARRYB_9__28_, CARRYB_9__27_,
         CARRYB_9__26_, CARRYB_9__25_, CARRYB_9__24_, CARRYB_9__23_,
         CARRYB_9__22_, CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_,
         CARRYB_9__18_, CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_,
         CARRYB_9__14_, CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_,
         CARRYB_9__10_, CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_,
         CARRYB_9__5_, CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_,
         CARRYB_9__0_, CARRYB_8__30_, CARRYB_8__29_, CARRYB_8__28_,
         CARRYB_8__27_, CARRYB_8__26_, CARRYB_8__25_, CARRYB_8__24_,
         CARRYB_8__23_, CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_,
         CARRYB_8__19_, CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_,
         CARRYB_8__15_, CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_,
         CARRYB_8__11_, CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_,
         CARRYB_8__7_, CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_,
         CARRYB_8__2_, CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__30_,
         CARRYB_7__29_, CARRYB_7__28_, CARRYB_7__27_, CARRYB_7__26_,
         CARRYB_7__25_, CARRYB_7__24_, CARRYB_7__23_, CARRYB_7__22_,
         CARRYB_7__21_, CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_,
         CARRYB_7__17_, CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_,
         CARRYB_7__13_, CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_,
         CARRYB_7__9_, CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_,
         CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_,
         CARRYB_6__30_, CARRYB_6__29_, CARRYB_6__28_, CARRYB_6__27_,
         CARRYB_6__26_, CARRYB_6__25_, CARRYB_6__24_, CARRYB_6__23_,
         CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_, CARRYB_6__19_,
         CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_, CARRYB_6__15_,
         CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_, CARRYB_6__11_,
         CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_, CARRYB_6__7_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__30_, CARRYB_5__29_, CARRYB_5__28_,
         CARRYB_5__27_, CARRYB_5__26_, CARRYB_5__25_, CARRYB_5__24_,
         CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_, CARRYB_5__20_,
         CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_, CARRYB_5__16_,
         CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_, CARRYB_5__12_,
         CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_, CARRYB_5__8_,
         CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__30_,
         CARRYB_4__29_, CARRYB_4__28_, CARRYB_4__27_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__30_, CARRYB_3__29_, CARRYB_3__28_, CARRYB_3__27_,
         CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_, CARRYB_3__23_,
         CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_, CARRYB_3__19_,
         CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_, CARRYB_3__15_,
         CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_, CARRYB_3__11_,
         CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_, CARRYB_3__7_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__30_, CARRYB_2__29_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_15__30_, SUMB_15__29_,
         SUMB_15__28_, SUMB_15__27_, SUMB_15__26_, SUMB_15__25_, SUMB_15__24_,
         SUMB_15__23_, SUMB_15__22_, SUMB_15__21_, SUMB_15__20_, SUMB_15__19_,
         SUMB_15__18_, SUMB_15__17_, SUMB_15__16_, SUMB_15__15_, SUMB_15__14_,
         SUMB_15__13_, SUMB_15__12_, SUMB_15__11_, SUMB_15__10_, SUMB_15__9_,
         SUMB_15__8_, SUMB_15__7_, SUMB_15__6_, SUMB_15__5_, SUMB_15__4_,
         SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__30_, SUMB_14__29_,
         SUMB_14__28_, SUMB_14__27_, SUMB_14__26_, SUMB_14__25_, SUMB_14__24_,
         SUMB_14__23_, SUMB_14__22_, SUMB_14__21_, SUMB_14__20_, SUMB_14__19_,
         SUMB_14__18_, SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_,
         SUMB_14__13_, SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_,
         SUMB_14__8_, SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_,
         SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__30_, SUMB_13__29_,
         SUMB_13__28_, SUMB_13__27_, SUMB_13__26_, SUMB_13__25_, SUMB_13__24_,
         SUMB_13__23_, SUMB_13__22_, SUMB_13__21_, SUMB_13__20_, SUMB_13__19_,
         SUMB_13__18_, SUMB_13__17_, SUMB_13__16_, SUMB_13__15_, SUMB_13__14_,
         SUMB_13__13_, SUMB_13__12_, SUMB_13__11_, SUMB_13__10_, SUMB_13__9_,
         SUMB_13__8_, SUMB_13__7_, SUMB_13__6_, SUMB_13__5_, SUMB_13__4_,
         SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__30_, SUMB_12__29_,
         SUMB_12__28_, SUMB_12__27_, SUMB_12__26_, SUMB_12__25_, SUMB_12__24_,
         SUMB_12__23_, SUMB_12__22_, SUMB_12__21_, SUMB_12__20_, SUMB_12__19_,
         SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_, SUMB_12__14_,
         SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_, SUMB_12__9_,
         SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_,
         SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__30_, SUMB_11__29_,
         SUMB_11__28_, SUMB_11__27_, SUMB_11__26_, SUMB_11__25_, SUMB_11__24_,
         SUMB_11__23_, SUMB_11__22_, SUMB_11__21_, SUMB_11__20_, SUMB_11__19_,
         SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_, SUMB_11__14_,
         SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_, SUMB_11__9_,
         SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__30_, SUMB_10__29_,
         SUMB_10__28_, SUMB_10__27_, SUMB_10__26_, SUMB_10__25_, SUMB_10__24_,
         SUMB_10__23_, SUMB_10__22_, SUMB_10__21_, SUMB_10__20_, SUMB_10__19_,
         SUMB_10__18_, SUMB_10__17_, SUMB_10__16_, SUMB_10__15_, SUMB_10__14_,
         SUMB_10__13_, SUMB_10__12_, SUMB_10__11_, SUMB_10__10_, SUMB_10__9_,
         SUMB_10__8_, SUMB_10__7_, SUMB_10__6_, SUMB_10__5_, SUMB_10__4_,
         SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__30_, SUMB_9__29_,
         SUMB_9__28_, SUMB_9__27_, SUMB_9__26_, SUMB_9__25_, SUMB_9__24_,
         SUMB_9__23_, SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_,
         SUMB_9__18_, SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_,
         SUMB_9__13_, SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_,
         SUMB_9__8_, SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_,
         SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__30_, SUMB_8__29_,
         SUMB_8__28_, SUMB_8__27_, SUMB_8__26_, SUMB_8__25_, SUMB_8__24_,
         SUMB_8__23_, SUMB_8__22_, SUMB_8__21_, SUMB_8__20_, SUMB_8__19_,
         SUMB_8__18_, SUMB_8__17_, SUMB_8__16_, SUMB_8__15_, SUMB_8__14_,
         SUMB_8__13_, SUMB_8__12_, SUMB_8__11_, SUMB_8__10_, SUMB_8__9_,
         SUMB_8__8_, SUMB_8__7_, SUMB_8__6_, SUMB_8__5_, SUMB_8__4_,
         SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__30_, SUMB_7__29_,
         SUMB_7__28_, SUMB_7__27_, SUMB_7__26_, SUMB_7__25_, SUMB_7__24_,
         SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_, SUMB_7__19_,
         SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_, SUMB_7__14_,
         SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_, SUMB_7__9_,
         SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_,
         SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__30_, SUMB_6__29_,
         SUMB_6__28_, SUMB_6__27_, SUMB_6__26_, SUMB_6__25_, SUMB_6__24_,
         SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_, SUMB_6__19_,
         SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_, SUMB_6__14_,
         SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_, SUMB_6__9_,
         SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__30_, SUMB_5__29_,
         SUMB_5__28_, SUMB_5__27_, SUMB_5__26_, SUMB_5__25_, SUMB_5__24_,
         SUMB_5__23_, SUMB_5__22_, SUMB_5__21_, SUMB_5__20_, SUMB_5__19_,
         SUMB_5__18_, SUMB_5__17_, SUMB_5__16_, SUMB_5__15_, SUMB_5__14_,
         SUMB_5__13_, SUMB_5__12_, SUMB_5__11_, SUMB_5__10_, SUMB_5__9_,
         SUMB_5__8_, SUMB_5__7_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__30_, SUMB_4__29_,
         SUMB_4__28_, SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_,
         SUMB_4__23_, SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_,
         SUMB_4__18_, SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_,
         SUMB_4__13_, SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_,
         SUMB_4__8_, SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_,
         SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__30_, SUMB_3__29_,
         SUMB_3__28_, SUMB_3__27_, SUMB_3__26_, SUMB_3__25_, SUMB_3__24_,
         SUMB_3__23_, SUMB_3__22_, SUMB_3__21_, SUMB_3__20_, SUMB_3__19_,
         SUMB_3__18_, SUMB_3__17_, SUMB_3__16_, SUMB_3__15_, SUMB_3__14_,
         SUMB_3__13_, SUMB_3__12_, SUMB_3__11_, SUMB_3__10_, SUMB_3__9_,
         SUMB_3__8_, SUMB_3__7_, SUMB_3__6_, SUMB_3__5_, SUMB_3__4_,
         SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__30_, SUMB_2__29_,
         SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_, SUMB_2__24_,
         SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_, SUMB_2__19_,
         SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_, SUMB_2__14_,
         SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_, SUMB_2__9_,
         SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_,
         SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, CARRYB_31__31_, CARRYB_31__30_,
         CARRYB_31__29_, CARRYB_31__28_, CARRYB_31__27_, CARRYB_31__26_,
         CARRYB_31__25_, CARRYB_31__24_, CARRYB_31__23_, CARRYB_31__22_,
         CARRYB_31__21_, CARRYB_31__20_, CARRYB_31__19_, CARRYB_31__18_,
         CARRYB_31__17_, CARRYB_31__16_, CARRYB_31__15_, CARRYB_31__14_,
         CARRYB_31__13_, CARRYB_31__12_, CARRYB_31__11_, CARRYB_31__10_,
         CARRYB_31__9_, CARRYB_31__8_, CARRYB_31__7_, CARRYB_31__6_,
         CARRYB_31__5_, CARRYB_31__4_, CARRYB_31__3_, CARRYB_31__2_,
         CARRYB_31__1_, CARRYB_31__0_, CARRYB_30__30_, CARRYB_30__29_,
         CARRYB_30__28_, CARRYB_30__27_, CARRYB_30__26_, CARRYB_30__25_,
         CARRYB_30__24_, CARRYB_30__23_, CARRYB_30__22_, CARRYB_30__21_,
         CARRYB_30__20_, CARRYB_30__19_, CARRYB_30__18_, CARRYB_30__17_,
         CARRYB_30__16_, CARRYB_30__15_, CARRYB_30__14_, CARRYB_30__13_,
         CARRYB_30__12_, CARRYB_30__11_, CARRYB_30__10_, CARRYB_30__9_,
         CARRYB_30__8_, CARRYB_30__7_, CARRYB_30__6_, CARRYB_30__5_,
         CARRYB_30__4_, CARRYB_30__3_, CARRYB_30__2_, CARRYB_30__1_,
         CARRYB_30__0_, CARRYB_29__30_, CARRYB_29__29_, CARRYB_29__28_,
         CARRYB_29__27_, CARRYB_29__26_, CARRYB_29__25_, CARRYB_29__24_,
         CARRYB_29__23_, CARRYB_29__22_, CARRYB_29__21_, CARRYB_29__20_,
         CARRYB_29__19_, CARRYB_29__18_, CARRYB_29__17_, CARRYB_29__16_,
         CARRYB_29__15_, CARRYB_29__14_, CARRYB_29__13_, CARRYB_29__12_,
         CARRYB_29__11_, CARRYB_29__10_, CARRYB_29__9_, CARRYB_29__8_,
         CARRYB_29__7_, CARRYB_29__6_, CARRYB_29__5_, CARRYB_29__4_,
         CARRYB_29__3_, CARRYB_29__2_, CARRYB_29__1_, CARRYB_29__0_,
         CARRYB_28__30_, CARRYB_28__29_, CARRYB_28__28_, CARRYB_28__27_,
         CARRYB_28__26_, CARRYB_28__25_, CARRYB_28__24_, CARRYB_28__23_,
         CARRYB_28__22_, CARRYB_28__21_, CARRYB_28__20_, CARRYB_28__19_,
         CARRYB_28__18_, CARRYB_28__17_, CARRYB_28__16_, CARRYB_28__15_,
         CARRYB_28__14_, CARRYB_28__13_, CARRYB_28__12_, CARRYB_28__11_,
         CARRYB_28__10_, CARRYB_28__9_, CARRYB_28__8_, CARRYB_28__7_,
         CARRYB_28__6_, CARRYB_28__5_, CARRYB_28__4_, CARRYB_28__3_,
         CARRYB_28__2_, CARRYB_28__1_, CARRYB_28__0_, CARRYB_27__30_,
         CARRYB_27__29_, CARRYB_27__28_, CARRYB_27__27_, CARRYB_27__26_,
         CARRYB_27__25_, CARRYB_27__24_, CARRYB_27__23_, CARRYB_27__22_,
         CARRYB_27__21_, CARRYB_27__20_, CARRYB_27__19_, CARRYB_27__18_,
         CARRYB_27__17_, CARRYB_27__16_, CARRYB_27__15_, CARRYB_27__14_,
         CARRYB_27__13_, CARRYB_27__12_, CARRYB_27__11_, CARRYB_27__10_,
         CARRYB_27__9_, CARRYB_27__8_, CARRYB_27__7_, CARRYB_27__6_,
         CARRYB_27__5_, CARRYB_27__4_, CARRYB_27__3_, CARRYB_27__2_,
         CARRYB_27__1_, CARRYB_27__0_, CARRYB_26__30_, CARRYB_26__29_,
         CARRYB_26__28_, CARRYB_26__27_, CARRYB_26__26_, CARRYB_26__25_,
         CARRYB_26__24_, CARRYB_26__23_, CARRYB_26__22_, CARRYB_26__21_,
         CARRYB_26__20_, CARRYB_26__19_, CARRYB_26__18_, CARRYB_26__17_,
         CARRYB_26__16_, CARRYB_26__15_, CARRYB_26__14_, CARRYB_26__13_,
         CARRYB_26__12_, CARRYB_26__11_, CARRYB_26__10_, CARRYB_26__9_,
         CARRYB_26__8_, CARRYB_26__7_, CARRYB_26__6_, CARRYB_26__5_,
         CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_, CARRYB_26__1_,
         CARRYB_26__0_, CARRYB_25__30_, CARRYB_25__29_, CARRYB_25__28_,
         CARRYB_25__27_, CARRYB_25__26_, CARRYB_25__25_, CARRYB_25__24_,
         CARRYB_25__23_, CARRYB_25__22_, CARRYB_25__21_, CARRYB_25__20_,
         CARRYB_25__19_, CARRYB_25__18_, CARRYB_25__17_, CARRYB_25__16_,
         CARRYB_25__15_, CARRYB_25__14_, CARRYB_25__13_, CARRYB_25__12_,
         CARRYB_25__11_, CARRYB_25__10_, CARRYB_25__9_, CARRYB_25__8_,
         CARRYB_25__7_, CARRYB_25__6_, CARRYB_25__5_, CARRYB_25__4_,
         CARRYB_25__3_, CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_,
         CARRYB_24__30_, CARRYB_24__29_, CARRYB_24__28_, CARRYB_24__27_,
         CARRYB_24__26_, CARRYB_24__25_, CARRYB_24__24_, CARRYB_24__23_,
         CARRYB_24__22_, CARRYB_24__21_, CARRYB_24__20_, CARRYB_24__19_,
         CARRYB_24__18_, CARRYB_24__17_, CARRYB_24__16_, CARRYB_24__15_,
         CARRYB_24__14_, CARRYB_24__13_, CARRYB_24__12_, CARRYB_24__11_,
         CARRYB_24__10_, CARRYB_24__9_, CARRYB_24__8_, CARRYB_24__7_,
         CARRYB_24__6_, CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_,
         CARRYB_24__2_, CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__30_,
         CARRYB_23__29_, CARRYB_23__28_, CARRYB_23__27_, CARRYB_23__26_,
         CARRYB_23__25_, CARRYB_23__24_, CARRYB_23__23_, CARRYB_23__22_,
         CARRYB_23__21_, CARRYB_23__20_, CARRYB_23__19_, CARRYB_23__18_,
         CARRYB_23__17_, CARRYB_23__16_, CARRYB_23__15_, CARRYB_23__14_,
         CARRYB_23__13_, CARRYB_23__12_, CARRYB_23__11_, CARRYB_23__10_,
         CARRYB_23__9_, CARRYB_23__8_, CARRYB_23__7_, CARRYB_23__6_,
         CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_, CARRYB_23__2_,
         CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__30_, CARRYB_22__29_,
         CARRYB_22__28_, CARRYB_22__27_, CARRYB_22__26_, CARRYB_22__25_,
         CARRYB_22__24_, CARRYB_22__23_, CARRYB_22__22_, CARRYB_22__21_,
         CARRYB_22__20_, CARRYB_22__19_, CARRYB_22__18_, CARRYB_22__17_,
         CARRYB_22__16_, CARRYB_22__15_, CARRYB_22__14_, CARRYB_22__13_,
         CARRYB_22__12_, CARRYB_22__11_, CARRYB_22__10_, CARRYB_22__9_,
         CARRYB_22__8_, CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_,
         CARRYB_22__4_, CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_,
         CARRYB_22__0_, CARRYB_21__30_, CARRYB_21__29_, CARRYB_21__28_,
         CARRYB_21__27_, CARRYB_21__26_, CARRYB_21__25_, CARRYB_21__24_,
         CARRYB_21__23_, CARRYB_21__22_, CARRYB_21__21_, CARRYB_21__20_,
         CARRYB_21__19_, CARRYB_21__18_, CARRYB_21__17_, CARRYB_21__16_,
         CARRYB_21__15_, CARRYB_21__14_, CARRYB_21__13_, CARRYB_21__12_,
         CARRYB_21__11_, CARRYB_21__10_, CARRYB_21__9_, CARRYB_21__8_,
         CARRYB_21__7_, CARRYB_21__6_, CARRYB_21__5_, CARRYB_21__4_,
         CARRYB_21__3_, CARRYB_21__2_, CARRYB_21__1_, CARRYB_21__0_,
         CARRYB_20__30_, CARRYB_20__29_, CARRYB_20__28_, CARRYB_20__27_,
         CARRYB_20__26_, CARRYB_20__25_, CARRYB_20__24_, CARRYB_20__23_,
         CARRYB_20__22_, CARRYB_20__21_, CARRYB_20__20_, CARRYB_20__19_,
         CARRYB_20__18_, CARRYB_20__17_, CARRYB_20__16_, CARRYB_20__15_,
         CARRYB_20__14_, CARRYB_20__13_, CARRYB_20__12_, CARRYB_20__11_,
         CARRYB_20__10_, CARRYB_20__9_, CARRYB_20__8_, CARRYB_20__7_,
         CARRYB_20__6_, CARRYB_20__5_, CARRYB_20__4_, CARRYB_20__3_,
         CARRYB_20__2_, CARRYB_20__1_, CARRYB_20__0_, CARRYB_19__30_,
         CARRYB_19__29_, CARRYB_19__28_, CARRYB_19__27_, CARRYB_19__26_,
         CARRYB_19__25_, CARRYB_19__24_, CARRYB_19__23_, CARRYB_19__22_,
         CARRYB_19__21_, CARRYB_19__20_, CARRYB_19__19_, CARRYB_19__18_,
         CARRYB_19__17_, CARRYB_19__16_, CARRYB_19__15_, CARRYB_19__14_,
         CARRYB_19__13_, CARRYB_19__12_, CARRYB_19__11_, CARRYB_19__10_,
         CARRYB_19__9_, CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_,
         CARRYB_19__5_, CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_,
         CARRYB_19__1_, CARRYB_19__0_, CARRYB_18__30_, CARRYB_18__29_,
         CARRYB_18__28_, CARRYB_18__27_, CARRYB_18__26_, CARRYB_18__25_,
         CARRYB_18__24_, CARRYB_18__23_, CARRYB_18__22_, CARRYB_18__21_,
         CARRYB_18__20_, CARRYB_18__19_, CARRYB_18__18_, CARRYB_18__17_,
         CARRYB_18__16_, CARRYB_18__15_, CARRYB_18__14_, CARRYB_18__13_,
         CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_, CARRYB_18__9_,
         CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_, CARRYB_18__5_,
         CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_, CARRYB_18__1_,
         CARRYB_18__0_, CARRYB_17__30_, CARRYB_17__29_, CARRYB_17__28_,
         CARRYB_17__27_, CARRYB_17__26_, CARRYB_17__25_, CARRYB_17__24_,
         CARRYB_17__23_, CARRYB_17__22_, CARRYB_17__21_, CARRYB_17__20_,
         CARRYB_17__19_, CARRYB_17__18_, CARRYB_17__17_, CARRYB_17__16_,
         CARRYB_17__15_, CARRYB_17__14_, CARRYB_17__13_, CARRYB_17__12_,
         CARRYB_17__11_, CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_,
         CARRYB_17__7_, CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_,
         CARRYB_17__3_, CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_,
         CARRYB_16__30_, CARRYB_16__29_, CARRYB_16__28_, CARRYB_16__27_,
         CARRYB_16__26_, CARRYB_16__25_, CARRYB_16__24_, CARRYB_16__23_,
         CARRYB_16__22_, CARRYB_16__21_, CARRYB_16__20_, CARRYB_16__19_,
         CARRYB_16__18_, CARRYB_16__17_, CARRYB_16__16_, CARRYB_16__15_,
         CARRYB_16__14_, CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_,
         CARRYB_16__10_, CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_,
         CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_,
         CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_, SUMB_31__31_,
         SUMB_31__30_, SUMB_31__29_, SUMB_31__28_, SUMB_31__27_, SUMB_31__26_,
         SUMB_31__25_, SUMB_31__24_, SUMB_31__23_, SUMB_31__22_, SUMB_31__21_,
         SUMB_31__20_, SUMB_31__19_, SUMB_31__18_, SUMB_31__17_, SUMB_31__16_,
         SUMB_31__15_, SUMB_31__14_, SUMB_31__13_, SUMB_31__12_, SUMB_31__11_,
         SUMB_31__10_, SUMB_31__9_, SUMB_31__8_, SUMB_31__7_, SUMB_31__6_,
         SUMB_31__5_, SUMB_31__4_, SUMB_31__3_, SUMB_31__2_, SUMB_31__1_,
         SUMB_31__0_, SUMB_30__30_, SUMB_30__29_, SUMB_30__28_, SUMB_30__27_,
         SUMB_30__26_, SUMB_30__25_, SUMB_30__24_, SUMB_30__23_, SUMB_30__22_,
         SUMB_30__21_, SUMB_30__20_, SUMB_30__19_, SUMB_30__18_, SUMB_30__17_,
         SUMB_30__16_, SUMB_30__15_, SUMB_30__14_, SUMB_30__13_, SUMB_30__12_,
         SUMB_30__11_, SUMB_30__10_, SUMB_30__9_, SUMB_30__8_, SUMB_30__7_,
         SUMB_30__6_, SUMB_30__5_, SUMB_30__4_, SUMB_30__3_, SUMB_30__2_,
         SUMB_30__1_, SUMB_29__30_, SUMB_29__29_, SUMB_29__28_, SUMB_29__27_,
         SUMB_29__26_, SUMB_29__25_, SUMB_29__24_, SUMB_29__23_, SUMB_29__22_,
         SUMB_29__21_, SUMB_29__20_, SUMB_29__19_, SUMB_29__18_, SUMB_29__17_,
         SUMB_29__16_, SUMB_29__15_, SUMB_29__14_, SUMB_29__13_, SUMB_29__12_,
         SUMB_29__11_, SUMB_29__10_, SUMB_29__9_, SUMB_29__8_, SUMB_29__7_,
         SUMB_29__6_, SUMB_29__5_, SUMB_29__4_, SUMB_29__3_, SUMB_29__2_,
         SUMB_29__1_, SUMB_28__30_, SUMB_28__29_, SUMB_28__28_, SUMB_28__27_,
         SUMB_28__26_, SUMB_28__25_, SUMB_28__24_, SUMB_28__23_, SUMB_28__22_,
         SUMB_28__21_, SUMB_28__20_, SUMB_28__19_, SUMB_28__18_, SUMB_28__17_,
         SUMB_28__16_, SUMB_28__15_, SUMB_28__14_, SUMB_28__13_, SUMB_28__12_,
         SUMB_28__11_, SUMB_28__10_, SUMB_28__9_, SUMB_28__8_, SUMB_28__7_,
         SUMB_28__6_, SUMB_28__5_, SUMB_28__4_, SUMB_28__3_, SUMB_28__2_,
         SUMB_28__1_, SUMB_27__30_, SUMB_27__29_, SUMB_27__28_, SUMB_27__27_,
         SUMB_27__26_, SUMB_27__25_, SUMB_27__24_, SUMB_27__23_, SUMB_27__22_,
         SUMB_27__21_, SUMB_27__20_, SUMB_27__19_, SUMB_27__18_, SUMB_27__17_,
         SUMB_27__16_, SUMB_27__15_, SUMB_27__14_, SUMB_27__13_, SUMB_27__12_,
         SUMB_27__11_, SUMB_27__10_, SUMB_27__9_, SUMB_27__8_, SUMB_27__7_,
         SUMB_27__6_, SUMB_27__5_, SUMB_27__4_, SUMB_27__3_, SUMB_27__2_,
         SUMB_27__1_, SUMB_26__30_, SUMB_26__29_, SUMB_26__28_, SUMB_26__27_,
         SUMB_26__26_, SUMB_26__25_, SUMB_26__24_, SUMB_26__23_, SUMB_26__22_,
         SUMB_26__21_, SUMB_26__20_, SUMB_26__19_, SUMB_26__18_, SUMB_26__17_,
         SUMB_26__16_, SUMB_26__15_, SUMB_26__14_, SUMB_26__13_, SUMB_26__12_,
         SUMB_26__11_, SUMB_26__10_, SUMB_26__9_, SUMB_26__8_, SUMB_26__7_,
         SUMB_26__6_, SUMB_26__5_, SUMB_26__4_, SUMB_26__3_, SUMB_26__2_,
         SUMB_26__1_, SUMB_25__30_, SUMB_25__29_, SUMB_25__28_, SUMB_25__27_,
         SUMB_25__26_, SUMB_25__25_, SUMB_25__24_, SUMB_25__23_, SUMB_25__22_,
         SUMB_25__21_, SUMB_25__20_, SUMB_25__19_, SUMB_25__18_, SUMB_25__17_,
         SUMB_25__16_, SUMB_25__15_, SUMB_25__14_, SUMB_25__13_, SUMB_25__12_,
         SUMB_25__11_, SUMB_25__10_, SUMB_25__9_, SUMB_25__8_, SUMB_25__7_,
         SUMB_25__6_, SUMB_25__5_, SUMB_25__4_, SUMB_25__3_, SUMB_25__2_,
         SUMB_25__1_, SUMB_24__30_, SUMB_24__29_, SUMB_24__28_, SUMB_24__27_,
         SUMB_24__26_, SUMB_24__25_, SUMB_24__24_, SUMB_24__23_, SUMB_24__22_,
         SUMB_24__21_, SUMB_24__20_, SUMB_24__19_, SUMB_24__18_, SUMB_24__17_,
         SUMB_24__16_, SUMB_24__15_, SUMB_24__14_, SUMB_24__13_, SUMB_24__12_,
         SUMB_24__11_, SUMB_24__10_, SUMB_24__9_, SUMB_24__8_, SUMB_24__7_,
         SUMB_24__6_, SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_,
         SUMB_24__1_, SUMB_23__30_, SUMB_23__29_, SUMB_23__28_, SUMB_23__27_,
         SUMB_23__26_, SUMB_23__25_, SUMB_23__24_, SUMB_23__23_, SUMB_23__22_,
         SUMB_23__21_, SUMB_23__20_, SUMB_23__19_, SUMB_23__18_, SUMB_23__17_,
         SUMB_23__16_, SUMB_23__15_, SUMB_23__14_, SUMB_23__13_, SUMB_23__12_,
         SUMB_23__11_, SUMB_23__10_, SUMB_23__9_, SUMB_23__8_, SUMB_23__7_,
         SUMB_23__6_, SUMB_23__5_, SUMB_23__4_, SUMB_23__3_, SUMB_23__2_,
         SUMB_23__1_, SUMB_22__30_, SUMB_22__29_, SUMB_22__28_, SUMB_22__27_,
         SUMB_22__26_, SUMB_22__25_, SUMB_22__24_, SUMB_22__23_, SUMB_22__22_,
         SUMB_22__21_, SUMB_22__20_, SUMB_22__19_, SUMB_22__18_, SUMB_22__17_,
         SUMB_22__16_, SUMB_22__15_, SUMB_22__14_, SUMB_22__13_, SUMB_22__12_,
         SUMB_22__11_, SUMB_22__10_, SUMB_22__9_, SUMB_22__8_, SUMB_22__7_,
         SUMB_22__6_, SUMB_22__5_, SUMB_22__4_, SUMB_22__3_, SUMB_22__2_,
         SUMB_22__1_, SUMB_21__30_, SUMB_21__29_, SUMB_21__28_, SUMB_21__27_,
         SUMB_21__26_, SUMB_21__25_, SUMB_21__24_, SUMB_21__23_, SUMB_21__22_,
         SUMB_21__21_, SUMB_21__20_, SUMB_21__19_, SUMB_21__18_, SUMB_21__17_,
         SUMB_21__16_, SUMB_21__15_, SUMB_21__14_, SUMB_21__13_, SUMB_21__12_,
         SUMB_21__11_, SUMB_21__10_, SUMB_21__9_, SUMB_21__8_, SUMB_21__7_,
         SUMB_21__6_, SUMB_21__5_, SUMB_21__4_, SUMB_21__3_, SUMB_21__2_,
         SUMB_21__1_, SUMB_20__30_, SUMB_20__29_, SUMB_20__28_, SUMB_20__27_,
         SUMB_20__26_, SUMB_20__25_, SUMB_20__24_, SUMB_20__23_, SUMB_20__22_,
         SUMB_20__21_, SUMB_20__20_, SUMB_20__19_, SUMB_20__18_, SUMB_20__17_,
         SUMB_20__16_, SUMB_20__15_, SUMB_20__14_, SUMB_20__13_, SUMB_20__12_,
         SUMB_20__11_, SUMB_20__10_, SUMB_20__9_, SUMB_20__8_, SUMB_20__7_,
         SUMB_20__6_, SUMB_20__5_, SUMB_20__4_, SUMB_20__3_, SUMB_20__2_,
         SUMB_20__1_, SUMB_19__30_, SUMB_19__29_, SUMB_19__28_, SUMB_19__27_,
         SUMB_19__26_, SUMB_19__25_, SUMB_19__24_, SUMB_19__23_, SUMB_19__22_,
         SUMB_19__21_, SUMB_19__20_, SUMB_19__19_, SUMB_19__18_, SUMB_19__17_,
         SUMB_19__16_, SUMB_19__15_, SUMB_19__14_, SUMB_19__13_, SUMB_19__12_,
         SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_,
         SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_,
         SUMB_19__1_, SUMB_18__30_, SUMB_18__29_, SUMB_18__28_, SUMB_18__27_,
         SUMB_18__26_, SUMB_18__25_, SUMB_18__24_, SUMB_18__23_, SUMB_18__22_,
         SUMB_18__21_, SUMB_18__20_, SUMB_18__19_, SUMB_18__18_, SUMB_18__17_,
         SUMB_18__16_, SUMB_18__15_, SUMB_18__14_, SUMB_18__13_, SUMB_18__12_,
         SUMB_18__11_, SUMB_18__10_, SUMB_18__9_, SUMB_18__8_, SUMB_18__7_,
         SUMB_18__6_, SUMB_18__5_, SUMB_18__4_, SUMB_18__3_, SUMB_18__2_,
         SUMB_18__1_, SUMB_17__30_, SUMB_17__29_, SUMB_17__28_, SUMB_17__27_,
         SUMB_17__26_, SUMB_17__25_, SUMB_17__24_, SUMB_17__23_, SUMB_17__22_,
         SUMB_17__21_, SUMB_17__20_, SUMB_17__19_, SUMB_17__18_, SUMB_17__17_,
         SUMB_17__16_, SUMB_17__15_, SUMB_17__14_, SUMB_17__13_, SUMB_17__12_,
         SUMB_17__11_, SUMB_17__10_, SUMB_17__9_, SUMB_17__8_, SUMB_17__7_,
         SUMB_17__6_, SUMB_17__5_, SUMB_17__4_, SUMB_17__3_, SUMB_17__2_,
         SUMB_17__1_, SUMB_16__30_, SUMB_16__29_, SUMB_16__28_, SUMB_16__27_,
         SUMB_16__26_, SUMB_16__25_, SUMB_16__24_, SUMB_16__23_, SUMB_16__22_,
         SUMB_16__21_, SUMB_16__20_, SUMB_16__19_, SUMB_16__18_, SUMB_16__17_,
         SUMB_16__16_, SUMB_16__15_, SUMB_16__14_, SUMB_16__13_, SUMB_16__12_,
         SUMB_16__11_, SUMB_16__10_, SUMB_16__9_, SUMB_16__8_, SUMB_16__7_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, A1_29_, A1_28_, A1_27_, A1_26_, A1_25_, A1_24_, A1_23_,
         A1_22_, A1_21_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_,
         A1_14_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_,
         A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_30_, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381;

  FA_X1 S14_31_0 ( .A(A[31]), .B(B[31]), .CI(SUMB_31__0_), .CO(A2_30_), .S(
        A1_29_) );
  FA_X1 S4_0 ( .A(ab_31__0_), .B(CARRYB_30__0_), .CI(SUMB_30__1_), .CO(
        CARRYB_31__0_), .S(SUMB_31__0_) );
  FA_X1 S4_1 ( .A(ab_31__1_), .B(CARRYB_30__1_), .CI(SUMB_30__2_), .CO(
        CARRYB_31__1_), .S(SUMB_31__1_) );
  FA_X1 S4_2 ( .A(ab_31__2_), .B(CARRYB_30__2_), .CI(SUMB_30__3_), .CO(
        CARRYB_31__2_), .S(SUMB_31__2_) );
  FA_X1 S4_3 ( .A(ab_31__3_), .B(CARRYB_30__3_), .CI(SUMB_30__4_), .CO(
        CARRYB_31__3_), .S(SUMB_31__3_) );
  FA_X1 S4_4 ( .A(ab_31__4_), .B(CARRYB_30__4_), .CI(SUMB_30__5_), .CO(
        CARRYB_31__4_), .S(SUMB_31__4_) );
  FA_X1 S4_5 ( .A(ab_31__5_), .B(CARRYB_30__5_), .CI(SUMB_30__6_), .CO(
        CARRYB_31__5_), .S(SUMB_31__5_) );
  FA_X1 S4_6 ( .A(ab_31__6_), .B(CARRYB_30__6_), .CI(SUMB_30__7_), .CO(
        CARRYB_31__6_), .S(SUMB_31__6_) );
  FA_X1 S4_7 ( .A(ab_31__7_), .B(CARRYB_30__7_), .CI(SUMB_30__8_), .CO(
        CARRYB_31__7_), .S(SUMB_31__7_) );
  FA_X1 S4_8 ( .A(ab_31__8_), .B(CARRYB_30__8_), .CI(SUMB_30__9_), .CO(
        CARRYB_31__8_), .S(SUMB_31__8_) );
  FA_X1 S4_9 ( .A(ab_31__9_), .B(CARRYB_30__9_), .CI(SUMB_30__10_), .CO(
        CARRYB_31__9_), .S(SUMB_31__9_) );
  FA_X1 S4_10 ( .A(ab_31__10_), .B(CARRYB_30__10_), .CI(SUMB_30__11_), .CO(
        CARRYB_31__10_), .S(SUMB_31__10_) );
  FA_X1 S4_11 ( .A(ab_31__11_), .B(CARRYB_30__11_), .CI(SUMB_30__12_), .CO(
        CARRYB_31__11_), .S(SUMB_31__11_) );
  FA_X1 S4_12 ( .A(ab_31__12_), .B(CARRYB_30__12_), .CI(SUMB_30__13_), .CO(
        CARRYB_31__12_), .S(SUMB_31__12_) );
  FA_X1 S4_13 ( .A(ab_31__13_), .B(CARRYB_30__13_), .CI(SUMB_30__14_), .CO(
        CARRYB_31__13_), .S(SUMB_31__13_) );
  FA_X1 S4_14 ( .A(ab_31__14_), .B(CARRYB_30__14_), .CI(SUMB_30__15_), .CO(
        CARRYB_31__14_), .S(SUMB_31__14_) );
  FA_X1 S4_15 ( .A(ab_31__15_), .B(CARRYB_30__15_), .CI(SUMB_30__16_), .CO(
        CARRYB_31__15_), .S(SUMB_31__15_) );
  FA_X1 S4_16 ( .A(ab_31__16_), .B(CARRYB_30__16_), .CI(SUMB_30__17_), .CO(
        CARRYB_31__16_), .S(SUMB_31__16_) );
  FA_X1 S4_17 ( .A(ab_31__17_), .B(CARRYB_30__17_), .CI(SUMB_30__18_), .CO(
        CARRYB_31__17_), .S(SUMB_31__17_) );
  FA_X1 S4_18 ( .A(ab_31__18_), .B(CARRYB_30__18_), .CI(SUMB_30__19_), .CO(
        CARRYB_31__18_), .S(SUMB_31__18_) );
  FA_X1 S4_19 ( .A(ab_31__19_), .B(CARRYB_30__19_), .CI(SUMB_30__20_), .CO(
        CARRYB_31__19_), .S(SUMB_31__19_) );
  FA_X1 S4_20 ( .A(ab_31__20_), .B(CARRYB_30__20_), .CI(SUMB_30__21_), .CO(
        CARRYB_31__20_), .S(SUMB_31__20_) );
  FA_X1 S4_21 ( .A(ab_31__21_), .B(CARRYB_30__21_), .CI(SUMB_30__22_), .CO(
        CARRYB_31__21_), .S(SUMB_31__21_) );
  FA_X1 S4_22 ( .A(ab_31__22_), .B(CARRYB_30__22_), .CI(SUMB_30__23_), .CO(
        CARRYB_31__22_), .S(SUMB_31__22_) );
  FA_X1 S4_23 ( .A(ab_31__23_), .B(CARRYB_30__23_), .CI(SUMB_30__24_), .CO(
        CARRYB_31__23_), .S(SUMB_31__23_) );
  FA_X1 S4_24 ( .A(ab_31__24_), .B(CARRYB_30__24_), .CI(SUMB_30__25_), .CO(
        CARRYB_31__24_), .S(SUMB_31__24_) );
  FA_X1 S4_25 ( .A(ab_31__25_), .B(CARRYB_30__25_), .CI(SUMB_30__26_), .CO(
        CARRYB_31__25_), .S(SUMB_31__25_) );
  FA_X1 S4_26 ( .A(ab_31__26_), .B(CARRYB_30__26_), .CI(SUMB_30__27_), .CO(
        CARRYB_31__26_), .S(SUMB_31__26_) );
  FA_X1 S4_27 ( .A(ab_31__27_), .B(CARRYB_30__27_), .CI(SUMB_30__28_), .CO(
        CARRYB_31__27_), .S(SUMB_31__27_) );
  FA_X1 S4_28 ( .A(ab_31__28_), .B(CARRYB_30__28_), .CI(SUMB_30__29_), .CO(
        CARRYB_31__28_), .S(SUMB_31__28_) );
  FA_X1 S4_29 ( .A(ab_31__29_), .B(CARRYB_30__29_), .CI(SUMB_30__30_), .CO(
        CARRYB_31__29_), .S(SUMB_31__29_) );
  FA_X1 S5_30 ( .A(ab_31__30_), .B(CARRYB_30__30_), .CI(ab_30__31_), .CO(
        CARRYB_31__30_), .S(SUMB_31__30_) );
  FA_X1 S14_31 ( .A(n222), .B(n127), .CI(ab_31__31_), .CO(CARRYB_31__31_), .S(
        SUMB_31__31_) );
  FA_X1 S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), .CO(
        CARRYB_30__0_), .S(A1_28_) );
  FA_X1 S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .CI(SUMB_29__2_), .CO(
        CARRYB_30__1_), .S(SUMB_30__1_) );
  FA_X1 S2_30_2 ( .A(ab_30__2_), .B(CARRYB_29__2_), .CI(SUMB_29__3_), .CO(
        CARRYB_30__2_), .S(SUMB_30__2_) );
  FA_X1 S2_30_3 ( .A(ab_30__3_), .B(CARRYB_29__3_), .CI(SUMB_29__4_), .CO(
        CARRYB_30__3_), .S(SUMB_30__3_) );
  FA_X1 S2_30_4 ( .A(ab_30__4_), .B(CARRYB_29__4_), .CI(SUMB_29__5_), .CO(
        CARRYB_30__4_), .S(SUMB_30__4_) );
  FA_X1 S2_30_5 ( .A(ab_30__5_), .B(CARRYB_29__5_), .CI(SUMB_29__6_), .CO(
        CARRYB_30__5_), .S(SUMB_30__5_) );
  FA_X1 S2_30_6 ( .A(ab_30__6_), .B(CARRYB_29__6_), .CI(SUMB_29__7_), .CO(
        CARRYB_30__6_), .S(SUMB_30__6_) );
  FA_X1 S2_30_7 ( .A(ab_30__7_), .B(CARRYB_29__7_), .CI(SUMB_29__8_), .CO(
        CARRYB_30__7_), .S(SUMB_30__7_) );
  FA_X1 S2_30_8 ( .A(ab_30__8_), .B(CARRYB_29__8_), .CI(SUMB_29__9_), .CO(
        CARRYB_30__8_), .S(SUMB_30__8_) );
  FA_X1 S2_30_9 ( .A(ab_30__9_), .B(CARRYB_29__9_), .CI(SUMB_29__10_), .CO(
        CARRYB_30__9_), .S(SUMB_30__9_) );
  FA_X1 S2_30_10 ( .A(ab_30__10_), .B(CARRYB_29__10_), .CI(SUMB_29__11_), .CO(
        CARRYB_30__10_), .S(SUMB_30__10_) );
  FA_X1 S2_30_11 ( .A(ab_30__11_), .B(CARRYB_29__11_), .CI(SUMB_29__12_), .CO(
        CARRYB_30__11_), .S(SUMB_30__11_) );
  FA_X1 S2_30_12 ( .A(ab_30__12_), .B(CARRYB_29__12_), .CI(SUMB_29__13_), .CO(
        CARRYB_30__12_), .S(SUMB_30__12_) );
  FA_X1 S2_30_13 ( .A(ab_30__13_), .B(CARRYB_29__13_), .CI(SUMB_29__14_), .CO(
        CARRYB_30__13_), .S(SUMB_30__13_) );
  FA_X1 S2_30_14 ( .A(ab_30__14_), .B(CARRYB_29__14_), .CI(SUMB_29__15_), .CO(
        CARRYB_30__14_), .S(SUMB_30__14_) );
  FA_X1 S2_30_15 ( .A(ab_30__15_), .B(CARRYB_29__15_), .CI(SUMB_29__16_), .CO(
        CARRYB_30__15_), .S(SUMB_30__15_) );
  FA_X1 S2_30_16 ( .A(ab_30__16_), .B(CARRYB_29__16_), .CI(SUMB_29__17_), .CO(
        CARRYB_30__16_), .S(SUMB_30__16_) );
  FA_X1 S2_30_17 ( .A(ab_30__17_), .B(CARRYB_29__17_), .CI(SUMB_29__18_), .CO(
        CARRYB_30__17_), .S(SUMB_30__17_) );
  FA_X1 S2_30_18 ( .A(ab_30__18_), .B(CARRYB_29__18_), .CI(SUMB_29__19_), .CO(
        CARRYB_30__18_), .S(SUMB_30__18_) );
  FA_X1 S2_30_19 ( .A(ab_30__19_), .B(CARRYB_29__19_), .CI(SUMB_29__20_), .CO(
        CARRYB_30__19_), .S(SUMB_30__19_) );
  FA_X1 S2_30_20 ( .A(ab_30__20_), .B(CARRYB_29__20_), .CI(SUMB_29__21_), .CO(
        CARRYB_30__20_), .S(SUMB_30__20_) );
  FA_X1 S2_30_21 ( .A(ab_30__21_), .B(CARRYB_29__21_), .CI(SUMB_29__22_), .CO(
        CARRYB_30__21_), .S(SUMB_30__21_) );
  FA_X1 S2_30_22 ( .A(ab_30__22_), .B(CARRYB_29__22_), .CI(SUMB_29__23_), .CO(
        CARRYB_30__22_), .S(SUMB_30__22_) );
  FA_X1 S2_30_23 ( .A(ab_30__23_), .B(CARRYB_29__23_), .CI(SUMB_29__24_), .CO(
        CARRYB_30__23_), .S(SUMB_30__23_) );
  FA_X1 S2_30_24 ( .A(ab_30__24_), .B(CARRYB_29__24_), .CI(SUMB_29__25_), .CO(
        CARRYB_30__24_), .S(SUMB_30__24_) );
  FA_X1 S2_30_25 ( .A(ab_30__25_), .B(CARRYB_29__25_), .CI(SUMB_29__26_), .CO(
        CARRYB_30__25_), .S(SUMB_30__25_) );
  FA_X1 S2_30_26 ( .A(ab_30__26_), .B(CARRYB_29__26_), .CI(SUMB_29__27_), .CO(
        CARRYB_30__26_), .S(SUMB_30__26_) );
  FA_X1 S2_30_27 ( .A(ab_30__27_), .B(CARRYB_29__27_), .CI(SUMB_29__28_), .CO(
        CARRYB_30__27_), .S(SUMB_30__27_) );
  FA_X1 S2_30_28 ( .A(ab_30__28_), .B(CARRYB_29__28_), .CI(SUMB_29__29_), .CO(
        CARRYB_30__28_), .S(SUMB_30__28_) );
  FA_X1 S2_30_29 ( .A(ab_30__29_), .B(CARRYB_29__29_), .CI(SUMB_29__30_), .CO(
        CARRYB_30__29_), .S(SUMB_30__29_) );
  FA_X1 S3_30_30 ( .A(ab_30__30_), .B(CARRYB_29__30_), .CI(ab_29__31_), .CO(
        CARRYB_30__30_), .S(SUMB_30__30_) );
  FA_X1 S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), .CO(
        CARRYB_29__0_), .S(A1_27_) );
  FA_X1 S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), .CO(
        CARRYB_29__1_), .S(SUMB_29__1_) );
  FA_X1 S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .CI(SUMB_28__3_), .CO(
        CARRYB_29__2_), .S(SUMB_29__2_) );
  FA_X1 S2_29_3 ( .A(ab_29__3_), .B(CARRYB_28__3_), .CI(SUMB_28__4_), .CO(
        CARRYB_29__3_), .S(SUMB_29__3_) );
  FA_X1 S2_29_4 ( .A(ab_29__4_), .B(CARRYB_28__4_), .CI(SUMB_28__5_), .CO(
        CARRYB_29__4_), .S(SUMB_29__4_) );
  FA_X1 S2_29_5 ( .A(ab_29__5_), .B(CARRYB_28__5_), .CI(SUMB_28__6_), .CO(
        CARRYB_29__5_), .S(SUMB_29__5_) );
  FA_X1 S2_29_6 ( .A(ab_29__6_), .B(CARRYB_28__6_), .CI(SUMB_28__7_), .CO(
        CARRYB_29__6_), .S(SUMB_29__6_) );
  FA_X1 S2_29_7 ( .A(ab_29__7_), .B(CARRYB_28__7_), .CI(SUMB_28__8_), .CO(
        CARRYB_29__7_), .S(SUMB_29__7_) );
  FA_X1 S2_29_8 ( .A(ab_29__8_), .B(CARRYB_28__8_), .CI(SUMB_28__9_), .CO(
        CARRYB_29__8_), .S(SUMB_29__8_) );
  FA_X1 S2_29_9 ( .A(ab_29__9_), .B(CARRYB_28__9_), .CI(SUMB_28__10_), .CO(
        CARRYB_29__9_), .S(SUMB_29__9_) );
  FA_X1 S2_29_10 ( .A(ab_29__10_), .B(CARRYB_28__10_), .CI(SUMB_28__11_), .CO(
        CARRYB_29__10_), .S(SUMB_29__10_) );
  FA_X1 S2_29_11 ( .A(ab_29__11_), .B(CARRYB_28__11_), .CI(SUMB_28__12_), .CO(
        CARRYB_29__11_), .S(SUMB_29__11_) );
  FA_X1 S2_29_12 ( .A(ab_29__12_), .B(CARRYB_28__12_), .CI(SUMB_28__13_), .CO(
        CARRYB_29__12_), .S(SUMB_29__12_) );
  FA_X1 S2_29_13 ( .A(ab_29__13_), .B(CARRYB_28__13_), .CI(SUMB_28__14_), .CO(
        CARRYB_29__13_), .S(SUMB_29__13_) );
  FA_X1 S2_29_14 ( .A(ab_29__14_), .B(CARRYB_28__14_), .CI(SUMB_28__15_), .CO(
        CARRYB_29__14_), .S(SUMB_29__14_) );
  FA_X1 S2_29_15 ( .A(ab_29__15_), .B(CARRYB_28__15_), .CI(SUMB_28__16_), .CO(
        CARRYB_29__15_), .S(SUMB_29__15_) );
  FA_X1 S2_29_16 ( .A(ab_29__16_), .B(CARRYB_28__16_), .CI(SUMB_28__17_), .CO(
        CARRYB_29__16_), .S(SUMB_29__16_) );
  FA_X1 S2_29_17 ( .A(ab_29__17_), .B(CARRYB_28__17_), .CI(SUMB_28__18_), .CO(
        CARRYB_29__17_), .S(SUMB_29__17_) );
  FA_X1 S2_29_18 ( .A(ab_29__18_), .B(CARRYB_28__18_), .CI(SUMB_28__19_), .CO(
        CARRYB_29__18_), .S(SUMB_29__18_) );
  FA_X1 S2_29_19 ( .A(ab_29__19_), .B(CARRYB_28__19_), .CI(SUMB_28__20_), .CO(
        CARRYB_29__19_), .S(SUMB_29__19_) );
  FA_X1 S2_29_20 ( .A(ab_29__20_), .B(CARRYB_28__20_), .CI(SUMB_28__21_), .CO(
        CARRYB_29__20_), .S(SUMB_29__20_) );
  FA_X1 S2_29_21 ( .A(ab_29__21_), .B(CARRYB_28__21_), .CI(SUMB_28__22_), .CO(
        CARRYB_29__21_), .S(SUMB_29__21_) );
  FA_X1 S2_29_22 ( .A(ab_29__22_), .B(CARRYB_28__22_), .CI(SUMB_28__23_), .CO(
        CARRYB_29__22_), .S(SUMB_29__22_) );
  FA_X1 S2_29_23 ( .A(ab_29__23_), .B(CARRYB_28__23_), .CI(SUMB_28__24_), .CO(
        CARRYB_29__23_), .S(SUMB_29__23_) );
  FA_X1 S2_29_24 ( .A(ab_29__24_), .B(CARRYB_28__24_), .CI(SUMB_28__25_), .CO(
        CARRYB_29__24_), .S(SUMB_29__24_) );
  FA_X1 S2_29_25 ( .A(ab_29__25_), .B(CARRYB_28__25_), .CI(SUMB_28__26_), .CO(
        CARRYB_29__25_), .S(SUMB_29__25_) );
  FA_X1 S2_29_26 ( .A(ab_29__26_), .B(CARRYB_28__26_), .CI(SUMB_28__27_), .CO(
        CARRYB_29__26_), .S(SUMB_29__26_) );
  FA_X1 S2_29_27 ( .A(ab_29__27_), .B(CARRYB_28__27_), .CI(SUMB_28__28_), .CO(
        CARRYB_29__27_), .S(SUMB_29__27_) );
  FA_X1 S2_29_28 ( .A(ab_29__28_), .B(CARRYB_28__28_), .CI(SUMB_28__29_), .CO(
        CARRYB_29__28_), .S(SUMB_29__28_) );
  FA_X1 S2_29_29 ( .A(ab_29__29_), .B(CARRYB_28__29_), .CI(SUMB_28__30_), .CO(
        CARRYB_29__29_), .S(SUMB_29__29_) );
  FA_X1 S3_29_30 ( .A(ab_29__30_), .B(CARRYB_28__30_), .CI(ab_28__31_), .CO(
        CARRYB_29__30_), .S(SUMB_29__30_) );
  FA_X1 S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), .CO(
        CARRYB_28__0_), .S(A1_26_) );
  FA_X1 S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), .CO(
        CARRYB_28__1_), .S(SUMB_28__1_) );
  FA_X1 S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), .CO(
        CARRYB_28__2_), .S(SUMB_28__2_) );
  FA_X1 S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .CI(SUMB_27__4_), .CO(
        CARRYB_28__3_), .S(SUMB_28__3_) );
  FA_X1 S2_28_4 ( .A(ab_28__4_), .B(CARRYB_27__4_), .CI(SUMB_27__5_), .CO(
        CARRYB_28__4_), .S(SUMB_28__4_) );
  FA_X1 S2_28_5 ( .A(ab_28__5_), .B(CARRYB_27__5_), .CI(SUMB_27__6_), .CO(
        CARRYB_28__5_), .S(SUMB_28__5_) );
  FA_X1 S2_28_6 ( .A(ab_28__6_), .B(CARRYB_27__6_), .CI(SUMB_27__7_), .CO(
        CARRYB_28__6_), .S(SUMB_28__6_) );
  FA_X1 S2_28_7 ( .A(ab_28__7_), .B(CARRYB_27__7_), .CI(SUMB_27__8_), .CO(
        CARRYB_28__7_), .S(SUMB_28__7_) );
  FA_X1 S2_28_8 ( .A(ab_28__8_), .B(CARRYB_27__8_), .CI(SUMB_27__9_), .CO(
        CARRYB_28__8_), .S(SUMB_28__8_) );
  FA_X1 S2_28_9 ( .A(ab_28__9_), .B(CARRYB_27__9_), .CI(SUMB_27__10_), .CO(
        CARRYB_28__9_), .S(SUMB_28__9_) );
  FA_X1 S2_28_10 ( .A(ab_28__10_), .B(CARRYB_27__10_), .CI(SUMB_27__11_), .CO(
        CARRYB_28__10_), .S(SUMB_28__10_) );
  FA_X1 S2_28_11 ( .A(ab_28__11_), .B(CARRYB_27__11_), .CI(SUMB_27__12_), .CO(
        CARRYB_28__11_), .S(SUMB_28__11_) );
  FA_X1 S2_28_12 ( .A(ab_28__12_), .B(CARRYB_27__12_), .CI(SUMB_27__13_), .CO(
        CARRYB_28__12_), .S(SUMB_28__12_) );
  FA_X1 S2_28_13 ( .A(ab_28__13_), .B(CARRYB_27__13_), .CI(SUMB_27__14_), .CO(
        CARRYB_28__13_), .S(SUMB_28__13_) );
  FA_X1 S2_28_14 ( .A(ab_28__14_), .B(CARRYB_27__14_), .CI(SUMB_27__15_), .CO(
        CARRYB_28__14_), .S(SUMB_28__14_) );
  FA_X1 S2_28_15 ( .A(ab_28__15_), .B(CARRYB_27__15_), .CI(SUMB_27__16_), .CO(
        CARRYB_28__15_), .S(SUMB_28__15_) );
  FA_X1 S2_28_16 ( .A(ab_28__16_), .B(CARRYB_27__16_), .CI(SUMB_27__17_), .CO(
        CARRYB_28__16_), .S(SUMB_28__16_) );
  FA_X1 S2_28_17 ( .A(ab_28__17_), .B(CARRYB_27__17_), .CI(SUMB_27__18_), .CO(
        CARRYB_28__17_), .S(SUMB_28__17_) );
  FA_X1 S2_28_18 ( .A(ab_28__18_), .B(CARRYB_27__18_), .CI(SUMB_27__19_), .CO(
        CARRYB_28__18_), .S(SUMB_28__18_) );
  FA_X1 S2_28_19 ( .A(ab_28__19_), .B(CARRYB_27__19_), .CI(SUMB_27__20_), .CO(
        CARRYB_28__19_), .S(SUMB_28__19_) );
  FA_X1 S2_28_20 ( .A(ab_28__20_), .B(CARRYB_27__20_), .CI(SUMB_27__21_), .CO(
        CARRYB_28__20_), .S(SUMB_28__20_) );
  FA_X1 S2_28_21 ( .A(ab_28__21_), .B(CARRYB_27__21_), .CI(SUMB_27__22_), .CO(
        CARRYB_28__21_), .S(SUMB_28__21_) );
  FA_X1 S2_28_22 ( .A(ab_28__22_), .B(CARRYB_27__22_), .CI(SUMB_27__23_), .CO(
        CARRYB_28__22_), .S(SUMB_28__22_) );
  FA_X1 S2_28_23 ( .A(ab_28__23_), .B(CARRYB_27__23_), .CI(SUMB_27__24_), .CO(
        CARRYB_28__23_), .S(SUMB_28__23_) );
  FA_X1 S2_28_24 ( .A(ab_28__24_), .B(CARRYB_27__24_), .CI(SUMB_27__25_), .CO(
        CARRYB_28__24_), .S(SUMB_28__24_) );
  FA_X1 S2_28_25 ( .A(ab_28__25_), .B(CARRYB_27__25_), .CI(SUMB_27__26_), .CO(
        CARRYB_28__25_), .S(SUMB_28__25_) );
  FA_X1 S2_28_26 ( .A(ab_28__26_), .B(CARRYB_27__26_), .CI(SUMB_27__27_), .CO(
        CARRYB_28__26_), .S(SUMB_28__26_) );
  FA_X1 S2_28_27 ( .A(ab_28__27_), .B(CARRYB_27__27_), .CI(SUMB_27__28_), .CO(
        CARRYB_28__27_), .S(SUMB_28__27_) );
  FA_X1 S2_28_28 ( .A(ab_28__28_), .B(CARRYB_27__28_), .CI(SUMB_27__29_), .CO(
        CARRYB_28__28_), .S(SUMB_28__28_) );
  FA_X1 S2_28_29 ( .A(ab_28__29_), .B(CARRYB_27__29_), .CI(SUMB_27__30_), .CO(
        CARRYB_28__29_), .S(SUMB_28__29_) );
  FA_X1 S3_28_30 ( .A(ab_28__30_), .B(CARRYB_27__30_), .CI(ab_27__31_), .CO(
        CARRYB_28__30_), .S(SUMB_28__30_) );
  FA_X1 S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), .CO(
        CARRYB_27__0_), .S(A1_25_) );
  FA_X1 S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), .CO(
        CARRYB_27__1_), .S(SUMB_27__1_) );
  FA_X1 S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), .CO(
        CARRYB_27__2_), .S(SUMB_27__2_) );
  FA_X1 S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), .CO(
        CARRYB_27__3_), .S(SUMB_27__3_) );
  FA_X1 S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .CI(SUMB_26__5_), .CO(
        CARRYB_27__4_), .S(SUMB_27__4_) );
  FA_X1 S2_27_5 ( .A(ab_27__5_), .B(CARRYB_26__5_), .CI(SUMB_26__6_), .CO(
        CARRYB_27__5_), .S(SUMB_27__5_) );
  FA_X1 S2_27_6 ( .A(ab_27__6_), .B(CARRYB_26__6_), .CI(SUMB_26__7_), .CO(
        CARRYB_27__6_), .S(SUMB_27__6_) );
  FA_X1 S2_27_7 ( .A(ab_27__7_), .B(CARRYB_26__7_), .CI(SUMB_26__8_), .CO(
        CARRYB_27__7_), .S(SUMB_27__7_) );
  FA_X1 S2_27_8 ( .A(ab_27__8_), .B(CARRYB_26__8_), .CI(SUMB_26__9_), .CO(
        CARRYB_27__8_), .S(SUMB_27__8_) );
  FA_X1 S2_27_9 ( .A(ab_27__9_), .B(CARRYB_26__9_), .CI(SUMB_26__10_), .CO(
        CARRYB_27__9_), .S(SUMB_27__9_) );
  FA_X1 S2_27_10 ( .A(ab_27__10_), .B(CARRYB_26__10_), .CI(SUMB_26__11_), .CO(
        CARRYB_27__10_), .S(SUMB_27__10_) );
  FA_X1 S2_27_11 ( .A(ab_27__11_), .B(CARRYB_26__11_), .CI(SUMB_26__12_), .CO(
        CARRYB_27__11_), .S(SUMB_27__11_) );
  FA_X1 S2_27_12 ( .A(ab_27__12_), .B(CARRYB_26__12_), .CI(SUMB_26__13_), .CO(
        CARRYB_27__12_), .S(SUMB_27__12_) );
  FA_X1 S2_27_13 ( .A(ab_27__13_), .B(CARRYB_26__13_), .CI(SUMB_26__14_), .CO(
        CARRYB_27__13_), .S(SUMB_27__13_) );
  FA_X1 S2_27_14 ( .A(ab_27__14_), .B(CARRYB_26__14_), .CI(SUMB_26__15_), .CO(
        CARRYB_27__14_), .S(SUMB_27__14_) );
  FA_X1 S2_27_15 ( .A(ab_27__15_), .B(CARRYB_26__15_), .CI(SUMB_26__16_), .CO(
        CARRYB_27__15_), .S(SUMB_27__15_) );
  FA_X1 S2_27_16 ( .A(ab_27__16_), .B(CARRYB_26__16_), .CI(SUMB_26__17_), .CO(
        CARRYB_27__16_), .S(SUMB_27__16_) );
  FA_X1 S2_27_17 ( .A(ab_27__17_), .B(CARRYB_26__17_), .CI(SUMB_26__18_), .CO(
        CARRYB_27__17_), .S(SUMB_27__17_) );
  FA_X1 S2_27_18 ( .A(ab_27__18_), .B(CARRYB_26__18_), .CI(SUMB_26__19_), .CO(
        CARRYB_27__18_), .S(SUMB_27__18_) );
  FA_X1 S2_27_19 ( .A(ab_27__19_), .B(CARRYB_26__19_), .CI(SUMB_26__20_), .CO(
        CARRYB_27__19_), .S(SUMB_27__19_) );
  FA_X1 S2_27_20 ( .A(ab_27__20_), .B(CARRYB_26__20_), .CI(SUMB_26__21_), .CO(
        CARRYB_27__20_), .S(SUMB_27__20_) );
  FA_X1 S2_27_21 ( .A(ab_27__21_), .B(CARRYB_26__21_), .CI(SUMB_26__22_), .CO(
        CARRYB_27__21_), .S(SUMB_27__21_) );
  FA_X1 S2_27_22 ( .A(ab_27__22_), .B(CARRYB_26__22_), .CI(SUMB_26__23_), .CO(
        CARRYB_27__22_), .S(SUMB_27__22_) );
  FA_X1 S2_27_23 ( .A(ab_27__23_), .B(CARRYB_26__23_), .CI(SUMB_26__24_), .CO(
        CARRYB_27__23_), .S(SUMB_27__23_) );
  FA_X1 S2_27_24 ( .A(ab_27__24_), .B(CARRYB_26__24_), .CI(SUMB_26__25_), .CO(
        CARRYB_27__24_), .S(SUMB_27__24_) );
  FA_X1 S2_27_25 ( .A(ab_27__25_), .B(CARRYB_26__25_), .CI(SUMB_26__26_), .CO(
        CARRYB_27__25_), .S(SUMB_27__25_) );
  FA_X1 S2_27_26 ( .A(ab_27__26_), .B(CARRYB_26__26_), .CI(SUMB_26__27_), .CO(
        CARRYB_27__26_), .S(SUMB_27__26_) );
  FA_X1 S2_27_27 ( .A(ab_27__27_), .B(CARRYB_26__27_), .CI(SUMB_26__28_), .CO(
        CARRYB_27__27_), .S(SUMB_27__27_) );
  FA_X1 S2_27_28 ( .A(ab_27__28_), .B(CARRYB_26__28_), .CI(SUMB_26__29_), .CO(
        CARRYB_27__28_), .S(SUMB_27__28_) );
  FA_X1 S2_27_29 ( .A(ab_27__29_), .B(CARRYB_26__29_), .CI(SUMB_26__30_), .CO(
        CARRYB_27__29_), .S(SUMB_27__29_) );
  FA_X1 S3_27_30 ( .A(ab_27__30_), .B(CARRYB_26__30_), .CI(ab_26__31_), .CO(
        CARRYB_27__30_), .S(SUMB_27__30_) );
  FA_X1 S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), .CO(
        CARRYB_26__0_), .S(A1_24_) );
  FA_X1 S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), .CO(
        CARRYB_26__1_), .S(SUMB_26__1_) );
  FA_X1 S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), .CO(
        CARRYB_26__2_), .S(SUMB_26__2_) );
  FA_X1 S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), .CO(
        CARRYB_26__3_), .S(SUMB_26__3_) );
  FA_X1 S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), .CO(
        CARRYB_26__4_), .S(SUMB_26__4_) );
  FA_X1 S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .CI(SUMB_25__6_), .CO(
        CARRYB_26__5_), .S(SUMB_26__5_) );
  FA_X1 S2_26_6 ( .A(ab_26__6_), .B(CARRYB_25__6_), .CI(SUMB_25__7_), .CO(
        CARRYB_26__6_), .S(SUMB_26__6_) );
  FA_X1 S2_26_7 ( .A(ab_26__7_), .B(CARRYB_25__7_), .CI(SUMB_25__8_), .CO(
        CARRYB_26__7_), .S(SUMB_26__7_) );
  FA_X1 S2_26_8 ( .A(ab_26__8_), .B(CARRYB_25__8_), .CI(SUMB_25__9_), .CO(
        CARRYB_26__8_), .S(SUMB_26__8_) );
  FA_X1 S2_26_9 ( .A(ab_26__9_), .B(CARRYB_25__9_), .CI(SUMB_25__10_), .CO(
        CARRYB_26__9_), .S(SUMB_26__9_) );
  FA_X1 S2_26_10 ( .A(ab_26__10_), .B(CARRYB_25__10_), .CI(SUMB_25__11_), .CO(
        CARRYB_26__10_), .S(SUMB_26__10_) );
  FA_X1 S2_26_11 ( .A(ab_26__11_), .B(CARRYB_25__11_), .CI(SUMB_25__12_), .CO(
        CARRYB_26__11_), .S(SUMB_26__11_) );
  FA_X1 S2_26_12 ( .A(ab_26__12_), .B(CARRYB_25__12_), .CI(SUMB_25__13_), .CO(
        CARRYB_26__12_), .S(SUMB_26__12_) );
  FA_X1 S2_26_13 ( .A(ab_26__13_), .B(CARRYB_25__13_), .CI(SUMB_25__14_), .CO(
        CARRYB_26__13_), .S(SUMB_26__13_) );
  FA_X1 S2_26_14 ( .A(ab_26__14_), .B(CARRYB_25__14_), .CI(SUMB_25__15_), .CO(
        CARRYB_26__14_), .S(SUMB_26__14_) );
  FA_X1 S2_26_15 ( .A(ab_26__15_), .B(CARRYB_25__15_), .CI(SUMB_25__16_), .CO(
        CARRYB_26__15_), .S(SUMB_26__15_) );
  FA_X1 S2_26_16 ( .A(ab_26__16_), .B(CARRYB_25__16_), .CI(SUMB_25__17_), .CO(
        CARRYB_26__16_), .S(SUMB_26__16_) );
  FA_X1 S2_26_17 ( .A(ab_26__17_), .B(CARRYB_25__17_), .CI(SUMB_25__18_), .CO(
        CARRYB_26__17_), .S(SUMB_26__17_) );
  FA_X1 S2_26_18 ( .A(ab_26__18_), .B(CARRYB_25__18_), .CI(SUMB_25__19_), .CO(
        CARRYB_26__18_), .S(SUMB_26__18_) );
  FA_X1 S2_26_19 ( .A(ab_26__19_), .B(CARRYB_25__19_), .CI(SUMB_25__20_), .CO(
        CARRYB_26__19_), .S(SUMB_26__19_) );
  FA_X1 S2_26_20 ( .A(ab_26__20_), .B(CARRYB_25__20_), .CI(SUMB_25__21_), .CO(
        CARRYB_26__20_), .S(SUMB_26__20_) );
  FA_X1 S2_26_21 ( .A(ab_26__21_), .B(CARRYB_25__21_), .CI(SUMB_25__22_), .CO(
        CARRYB_26__21_), .S(SUMB_26__21_) );
  FA_X1 S2_26_22 ( .A(ab_26__22_), .B(CARRYB_25__22_), .CI(SUMB_25__23_), .CO(
        CARRYB_26__22_), .S(SUMB_26__22_) );
  FA_X1 S2_26_23 ( .A(ab_26__23_), .B(CARRYB_25__23_), .CI(SUMB_25__24_), .CO(
        CARRYB_26__23_), .S(SUMB_26__23_) );
  FA_X1 S2_26_24 ( .A(ab_26__24_), .B(CARRYB_25__24_), .CI(SUMB_25__25_), .CO(
        CARRYB_26__24_), .S(SUMB_26__24_) );
  FA_X1 S2_26_25 ( .A(ab_26__25_), .B(CARRYB_25__25_), .CI(SUMB_25__26_), .CO(
        CARRYB_26__25_), .S(SUMB_26__25_) );
  FA_X1 S2_26_26 ( .A(ab_26__26_), .B(CARRYB_25__26_), .CI(SUMB_25__27_), .CO(
        CARRYB_26__26_), .S(SUMB_26__26_) );
  FA_X1 S2_26_27 ( .A(ab_26__27_), .B(CARRYB_25__27_), .CI(SUMB_25__28_), .CO(
        CARRYB_26__27_), .S(SUMB_26__27_) );
  FA_X1 S2_26_28 ( .A(ab_26__28_), .B(CARRYB_25__28_), .CI(SUMB_25__29_), .CO(
        CARRYB_26__28_), .S(SUMB_26__28_) );
  FA_X1 S2_26_29 ( .A(ab_26__29_), .B(CARRYB_25__29_), .CI(SUMB_25__30_), .CO(
        CARRYB_26__29_), .S(SUMB_26__29_) );
  FA_X1 S3_26_30 ( .A(ab_26__30_), .B(CARRYB_25__30_), .CI(ab_25__31_), .CO(
        CARRYB_26__30_), .S(SUMB_26__30_) );
  FA_X1 S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), .CO(
        CARRYB_25__0_), .S(A1_23_) );
  FA_X1 S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), .CO(
        CARRYB_25__1_), .S(SUMB_25__1_) );
  FA_X1 S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), .CO(
        CARRYB_25__2_), .S(SUMB_25__2_) );
  FA_X1 S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), .CO(
        CARRYB_25__3_), .S(SUMB_25__3_) );
  FA_X1 S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), .CO(
        CARRYB_25__4_), .S(SUMB_25__4_) );
  FA_X1 S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), .CO(
        CARRYB_25__5_), .S(SUMB_25__5_) );
  FA_X1 S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .CI(SUMB_24__7_), .CO(
        CARRYB_25__6_), .S(SUMB_25__6_) );
  FA_X1 S2_25_7 ( .A(ab_25__7_), .B(CARRYB_24__7_), .CI(SUMB_24__8_), .CO(
        CARRYB_25__7_), .S(SUMB_25__7_) );
  FA_X1 S2_25_8 ( .A(ab_25__8_), .B(CARRYB_24__8_), .CI(SUMB_24__9_), .CO(
        CARRYB_25__8_), .S(SUMB_25__8_) );
  FA_X1 S2_25_9 ( .A(ab_25__9_), .B(CARRYB_24__9_), .CI(SUMB_24__10_), .CO(
        CARRYB_25__9_), .S(SUMB_25__9_) );
  FA_X1 S2_25_10 ( .A(ab_25__10_), .B(CARRYB_24__10_), .CI(SUMB_24__11_), .CO(
        CARRYB_25__10_), .S(SUMB_25__10_) );
  FA_X1 S2_25_11 ( .A(ab_25__11_), .B(CARRYB_24__11_), .CI(SUMB_24__12_), .CO(
        CARRYB_25__11_), .S(SUMB_25__11_) );
  FA_X1 S2_25_12 ( .A(ab_25__12_), .B(CARRYB_24__12_), .CI(SUMB_24__13_), .CO(
        CARRYB_25__12_), .S(SUMB_25__12_) );
  FA_X1 S2_25_13 ( .A(ab_25__13_), .B(CARRYB_24__13_), .CI(SUMB_24__14_), .CO(
        CARRYB_25__13_), .S(SUMB_25__13_) );
  FA_X1 S2_25_14 ( .A(ab_25__14_), .B(CARRYB_24__14_), .CI(SUMB_24__15_), .CO(
        CARRYB_25__14_), .S(SUMB_25__14_) );
  FA_X1 S2_25_15 ( .A(ab_25__15_), .B(CARRYB_24__15_), .CI(SUMB_24__16_), .CO(
        CARRYB_25__15_), .S(SUMB_25__15_) );
  FA_X1 S2_25_16 ( .A(ab_25__16_), .B(CARRYB_24__16_), .CI(SUMB_24__17_), .CO(
        CARRYB_25__16_), .S(SUMB_25__16_) );
  FA_X1 S2_25_17 ( .A(ab_25__17_), .B(CARRYB_24__17_), .CI(SUMB_24__18_), .CO(
        CARRYB_25__17_), .S(SUMB_25__17_) );
  FA_X1 S2_25_18 ( .A(ab_25__18_), .B(CARRYB_24__18_), .CI(SUMB_24__19_), .CO(
        CARRYB_25__18_), .S(SUMB_25__18_) );
  FA_X1 S2_25_19 ( .A(ab_25__19_), .B(CARRYB_24__19_), .CI(SUMB_24__20_), .CO(
        CARRYB_25__19_), .S(SUMB_25__19_) );
  FA_X1 S2_25_20 ( .A(ab_25__20_), .B(CARRYB_24__20_), .CI(SUMB_24__21_), .CO(
        CARRYB_25__20_), .S(SUMB_25__20_) );
  FA_X1 S2_25_21 ( .A(ab_25__21_), .B(CARRYB_24__21_), .CI(SUMB_24__22_), .CO(
        CARRYB_25__21_), .S(SUMB_25__21_) );
  FA_X1 S2_25_22 ( .A(ab_25__22_), .B(CARRYB_24__22_), .CI(SUMB_24__23_), .CO(
        CARRYB_25__22_), .S(SUMB_25__22_) );
  FA_X1 S2_25_23 ( .A(ab_25__23_), .B(CARRYB_24__23_), .CI(SUMB_24__24_), .CO(
        CARRYB_25__23_), .S(SUMB_25__23_) );
  FA_X1 S2_25_24 ( .A(ab_25__24_), .B(CARRYB_24__24_), .CI(SUMB_24__25_), .CO(
        CARRYB_25__24_), .S(SUMB_25__24_) );
  FA_X1 S2_25_25 ( .A(ab_25__25_), .B(CARRYB_24__25_), .CI(SUMB_24__26_), .CO(
        CARRYB_25__25_), .S(SUMB_25__25_) );
  FA_X1 S2_25_26 ( .A(ab_25__26_), .B(CARRYB_24__26_), .CI(SUMB_24__27_), .CO(
        CARRYB_25__26_), .S(SUMB_25__26_) );
  FA_X1 S2_25_27 ( .A(ab_25__27_), .B(CARRYB_24__27_), .CI(SUMB_24__28_), .CO(
        CARRYB_25__27_), .S(SUMB_25__27_) );
  FA_X1 S2_25_28 ( .A(ab_25__28_), .B(CARRYB_24__28_), .CI(SUMB_24__29_), .CO(
        CARRYB_25__28_), .S(SUMB_25__28_) );
  FA_X1 S2_25_29 ( .A(ab_25__29_), .B(CARRYB_24__29_), .CI(SUMB_24__30_), .CO(
        CARRYB_25__29_), .S(SUMB_25__29_) );
  FA_X1 S3_25_30 ( .A(ab_25__30_), .B(CARRYB_24__30_), .CI(ab_24__31_), .CO(
        CARRYB_25__30_), .S(SUMB_25__30_) );
  FA_X1 S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), .CO(
        CARRYB_24__0_), .S(A1_22_) );
  FA_X1 S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), .CO(
        CARRYB_24__1_), .S(SUMB_24__1_) );
  FA_X1 S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), .CO(
        CARRYB_24__2_), .S(SUMB_24__2_) );
  FA_X1 S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), .CO(
        CARRYB_24__3_), .S(SUMB_24__3_) );
  FA_X1 S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), .CO(
        CARRYB_24__4_), .S(SUMB_24__4_) );
  FA_X1 S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), .CO(
        CARRYB_24__5_), .S(SUMB_24__5_) );
  FA_X1 S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), .CO(
        CARRYB_24__6_), .S(SUMB_24__6_) );
  FA_X1 S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .CI(SUMB_23__8_), .CO(
        CARRYB_24__7_), .S(SUMB_24__7_) );
  FA_X1 S2_24_8 ( .A(ab_24__8_), .B(CARRYB_23__8_), .CI(SUMB_23__9_), .CO(
        CARRYB_24__8_), .S(SUMB_24__8_) );
  FA_X1 S2_24_9 ( .A(ab_24__9_), .B(CARRYB_23__9_), .CI(SUMB_23__10_), .CO(
        CARRYB_24__9_), .S(SUMB_24__9_) );
  FA_X1 S2_24_10 ( .A(ab_24__10_), .B(CARRYB_23__10_), .CI(SUMB_23__11_), .CO(
        CARRYB_24__10_), .S(SUMB_24__10_) );
  FA_X1 S2_24_11 ( .A(ab_24__11_), .B(CARRYB_23__11_), .CI(SUMB_23__12_), .CO(
        CARRYB_24__11_), .S(SUMB_24__11_) );
  FA_X1 S2_24_12 ( .A(ab_24__12_), .B(CARRYB_23__12_), .CI(SUMB_23__13_), .CO(
        CARRYB_24__12_), .S(SUMB_24__12_) );
  FA_X1 S2_24_13 ( .A(ab_24__13_), .B(CARRYB_23__13_), .CI(SUMB_23__14_), .CO(
        CARRYB_24__13_), .S(SUMB_24__13_) );
  FA_X1 S2_24_14 ( .A(ab_24__14_), .B(CARRYB_23__14_), .CI(SUMB_23__15_), .CO(
        CARRYB_24__14_), .S(SUMB_24__14_) );
  FA_X1 S2_24_15 ( .A(ab_24__15_), .B(CARRYB_23__15_), .CI(SUMB_23__16_), .CO(
        CARRYB_24__15_), .S(SUMB_24__15_) );
  FA_X1 S2_24_16 ( .A(ab_24__16_), .B(CARRYB_23__16_), .CI(SUMB_23__17_), .CO(
        CARRYB_24__16_), .S(SUMB_24__16_) );
  FA_X1 S2_24_17 ( .A(ab_24__17_), .B(CARRYB_23__17_), .CI(SUMB_23__18_), .CO(
        CARRYB_24__17_), .S(SUMB_24__17_) );
  FA_X1 S2_24_18 ( .A(ab_24__18_), .B(CARRYB_23__18_), .CI(SUMB_23__19_), .CO(
        CARRYB_24__18_), .S(SUMB_24__18_) );
  FA_X1 S2_24_19 ( .A(ab_24__19_), .B(CARRYB_23__19_), .CI(SUMB_23__20_), .CO(
        CARRYB_24__19_), .S(SUMB_24__19_) );
  FA_X1 S2_24_20 ( .A(ab_24__20_), .B(CARRYB_23__20_), .CI(SUMB_23__21_), .CO(
        CARRYB_24__20_), .S(SUMB_24__20_) );
  FA_X1 S2_24_21 ( .A(ab_24__21_), .B(CARRYB_23__21_), .CI(SUMB_23__22_), .CO(
        CARRYB_24__21_), .S(SUMB_24__21_) );
  FA_X1 S2_24_22 ( .A(ab_24__22_), .B(CARRYB_23__22_), .CI(SUMB_23__23_), .CO(
        CARRYB_24__22_), .S(SUMB_24__22_) );
  FA_X1 S2_24_23 ( .A(ab_24__23_), .B(CARRYB_23__23_), .CI(SUMB_23__24_), .CO(
        CARRYB_24__23_), .S(SUMB_24__23_) );
  FA_X1 S2_24_24 ( .A(ab_24__24_), .B(CARRYB_23__24_), .CI(SUMB_23__25_), .CO(
        CARRYB_24__24_), .S(SUMB_24__24_) );
  FA_X1 S2_24_25 ( .A(ab_24__25_), .B(CARRYB_23__25_), .CI(SUMB_23__26_), .CO(
        CARRYB_24__25_), .S(SUMB_24__25_) );
  FA_X1 S2_24_26 ( .A(ab_24__26_), .B(CARRYB_23__26_), .CI(SUMB_23__27_), .CO(
        CARRYB_24__26_), .S(SUMB_24__26_) );
  FA_X1 S2_24_27 ( .A(ab_24__27_), .B(CARRYB_23__27_), .CI(SUMB_23__28_), .CO(
        CARRYB_24__27_), .S(SUMB_24__27_) );
  FA_X1 S2_24_28 ( .A(ab_24__28_), .B(CARRYB_23__28_), .CI(SUMB_23__29_), .CO(
        CARRYB_24__28_), .S(SUMB_24__28_) );
  FA_X1 S2_24_29 ( .A(ab_24__29_), .B(CARRYB_23__29_), .CI(SUMB_23__30_), .CO(
        CARRYB_24__29_), .S(SUMB_24__29_) );
  FA_X1 S3_24_30 ( .A(ab_24__30_), .B(CARRYB_23__30_), .CI(ab_23__31_), .CO(
        CARRYB_24__30_), .S(SUMB_24__30_) );
  FA_X1 S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), .CO(
        CARRYB_23__0_), .S(A1_21_) );
  FA_X1 S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), .CO(
        CARRYB_23__1_), .S(SUMB_23__1_) );
  FA_X1 S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), .CO(
        CARRYB_23__2_), .S(SUMB_23__2_) );
  FA_X1 S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), .CO(
        CARRYB_23__3_), .S(SUMB_23__3_) );
  FA_X1 S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), .CO(
        CARRYB_23__4_), .S(SUMB_23__4_) );
  FA_X1 S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), .CO(
        CARRYB_23__5_), .S(SUMB_23__5_) );
  FA_X1 S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), .CO(
        CARRYB_23__6_), .S(SUMB_23__6_) );
  FA_X1 S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), .CO(
        CARRYB_23__7_), .S(SUMB_23__7_) );
  FA_X1 S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .CO(
        CARRYB_23__8_), .S(SUMB_23__8_) );
  FA_X1 S2_23_9 ( .A(ab_23__9_), .B(CARRYB_22__9_), .CI(SUMB_22__10_), .CO(
        CARRYB_23__9_), .S(SUMB_23__9_) );
  FA_X1 S2_23_10 ( .A(ab_23__10_), .B(CARRYB_22__10_), .CI(SUMB_22__11_), .CO(
        CARRYB_23__10_), .S(SUMB_23__10_) );
  FA_X1 S2_23_11 ( .A(ab_23__11_), .B(CARRYB_22__11_), .CI(SUMB_22__12_), .CO(
        CARRYB_23__11_), .S(SUMB_23__11_) );
  FA_X1 S2_23_12 ( .A(ab_23__12_), .B(CARRYB_22__12_), .CI(SUMB_22__13_), .CO(
        CARRYB_23__12_), .S(SUMB_23__12_) );
  FA_X1 S2_23_13 ( .A(ab_23__13_), .B(CARRYB_22__13_), .CI(SUMB_22__14_), .CO(
        CARRYB_23__13_), .S(SUMB_23__13_) );
  FA_X1 S2_23_14 ( .A(ab_23__14_), .B(CARRYB_22__14_), .CI(SUMB_22__15_), .CO(
        CARRYB_23__14_), .S(SUMB_23__14_) );
  FA_X1 S2_23_15 ( .A(ab_23__15_), .B(CARRYB_22__15_), .CI(SUMB_22__16_), .CO(
        CARRYB_23__15_), .S(SUMB_23__15_) );
  FA_X1 S2_23_16 ( .A(ab_23__16_), .B(CARRYB_22__16_), .CI(SUMB_22__17_), .CO(
        CARRYB_23__16_), .S(SUMB_23__16_) );
  FA_X1 S2_23_17 ( .A(ab_23__17_), .B(CARRYB_22__17_), .CI(SUMB_22__18_), .CO(
        CARRYB_23__17_), .S(SUMB_23__17_) );
  FA_X1 S2_23_18 ( .A(ab_23__18_), .B(CARRYB_22__18_), .CI(SUMB_22__19_), .CO(
        CARRYB_23__18_), .S(SUMB_23__18_) );
  FA_X1 S2_23_19 ( .A(ab_23__19_), .B(CARRYB_22__19_), .CI(SUMB_22__20_), .CO(
        CARRYB_23__19_), .S(SUMB_23__19_) );
  FA_X1 S2_23_20 ( .A(ab_23__20_), .B(CARRYB_22__20_), .CI(SUMB_22__21_), .CO(
        CARRYB_23__20_), .S(SUMB_23__20_) );
  FA_X1 S2_23_21 ( .A(ab_23__21_), .B(CARRYB_22__21_), .CI(SUMB_22__22_), .CO(
        CARRYB_23__21_), .S(SUMB_23__21_) );
  FA_X1 S2_23_22 ( .A(ab_23__22_), .B(CARRYB_22__22_), .CI(SUMB_22__23_), .CO(
        CARRYB_23__22_), .S(SUMB_23__22_) );
  FA_X1 S2_23_23 ( .A(ab_23__23_), .B(CARRYB_22__23_), .CI(SUMB_22__24_), .CO(
        CARRYB_23__23_), .S(SUMB_23__23_) );
  FA_X1 S2_23_24 ( .A(ab_23__24_), .B(CARRYB_22__24_), .CI(SUMB_22__25_), .CO(
        CARRYB_23__24_), .S(SUMB_23__24_) );
  FA_X1 S2_23_25 ( .A(ab_23__25_), .B(CARRYB_22__25_), .CI(SUMB_22__26_), .CO(
        CARRYB_23__25_), .S(SUMB_23__25_) );
  FA_X1 S2_23_26 ( .A(ab_23__26_), .B(CARRYB_22__26_), .CI(SUMB_22__27_), .CO(
        CARRYB_23__26_), .S(SUMB_23__26_) );
  FA_X1 S2_23_27 ( .A(ab_23__27_), .B(CARRYB_22__27_), .CI(SUMB_22__28_), .CO(
        CARRYB_23__27_), .S(SUMB_23__27_) );
  FA_X1 S2_23_28 ( .A(ab_23__28_), .B(CARRYB_22__28_), .CI(SUMB_22__29_), .CO(
        CARRYB_23__28_), .S(SUMB_23__28_) );
  FA_X1 S2_23_29 ( .A(ab_23__29_), .B(CARRYB_22__29_), .CI(SUMB_22__30_), .CO(
        CARRYB_23__29_), .S(SUMB_23__29_) );
  FA_X1 S3_23_30 ( .A(ab_23__30_), .B(CARRYB_22__30_), .CI(ab_22__31_), .CO(
        CARRYB_23__30_), .S(SUMB_23__30_) );
  FA_X1 S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), .CO(
        CARRYB_22__0_), .S(A1_20_) );
  FA_X1 S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), .CO(
        CARRYB_22__1_), .S(SUMB_22__1_) );
  FA_X1 S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), .CO(
        CARRYB_22__2_), .S(SUMB_22__2_) );
  FA_X1 S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), .CO(
        CARRYB_22__3_), .S(SUMB_22__3_) );
  FA_X1 S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), .CO(
        CARRYB_22__4_), .S(SUMB_22__4_) );
  FA_X1 S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), .CO(
        CARRYB_22__5_), .S(SUMB_22__5_) );
  FA_X1 S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), .CO(
        CARRYB_22__6_), .S(SUMB_22__6_) );
  FA_X1 S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), .CO(
        CARRYB_22__7_), .S(SUMB_22__7_) );
  FA_X1 S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), .CO(
        CARRYB_22__8_), .S(SUMB_22__8_) );
  FA_X1 S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), .CO(
        CARRYB_22__9_), .S(SUMB_22__9_) );
  FA_X1 S2_22_10 ( .A(ab_22__10_), .B(CARRYB_21__10_), .CI(SUMB_21__11_), .CO(
        CARRYB_22__10_), .S(SUMB_22__10_) );
  FA_X1 S2_22_11 ( .A(ab_22__11_), .B(CARRYB_21__11_), .CI(SUMB_21__12_), .CO(
        CARRYB_22__11_), .S(SUMB_22__11_) );
  FA_X1 S2_22_12 ( .A(ab_22__12_), .B(CARRYB_21__12_), .CI(SUMB_21__13_), .CO(
        CARRYB_22__12_), .S(SUMB_22__12_) );
  FA_X1 S2_22_13 ( .A(ab_22__13_), .B(CARRYB_21__13_), .CI(SUMB_21__14_), .CO(
        CARRYB_22__13_), .S(SUMB_22__13_) );
  FA_X1 S2_22_14 ( .A(ab_22__14_), .B(CARRYB_21__14_), .CI(SUMB_21__15_), .CO(
        CARRYB_22__14_), .S(SUMB_22__14_) );
  FA_X1 S2_22_15 ( .A(ab_22__15_), .B(CARRYB_21__15_), .CI(SUMB_21__16_), .CO(
        CARRYB_22__15_), .S(SUMB_22__15_) );
  FA_X1 S2_22_16 ( .A(ab_22__16_), .B(CARRYB_21__16_), .CI(SUMB_21__17_), .CO(
        CARRYB_22__16_), .S(SUMB_22__16_) );
  FA_X1 S2_22_17 ( .A(ab_22__17_), .B(CARRYB_21__17_), .CI(SUMB_21__18_), .CO(
        CARRYB_22__17_), .S(SUMB_22__17_) );
  FA_X1 S2_22_18 ( .A(ab_22__18_), .B(CARRYB_21__18_), .CI(SUMB_21__19_), .CO(
        CARRYB_22__18_), .S(SUMB_22__18_) );
  FA_X1 S2_22_19 ( .A(ab_22__19_), .B(CARRYB_21__19_), .CI(SUMB_21__20_), .CO(
        CARRYB_22__19_), .S(SUMB_22__19_) );
  FA_X1 S2_22_20 ( .A(ab_22__20_), .B(CARRYB_21__20_), .CI(SUMB_21__21_), .CO(
        CARRYB_22__20_), .S(SUMB_22__20_) );
  FA_X1 S2_22_21 ( .A(ab_22__21_), .B(CARRYB_21__21_), .CI(SUMB_21__22_), .CO(
        CARRYB_22__21_), .S(SUMB_22__21_) );
  FA_X1 S2_22_22 ( .A(ab_22__22_), .B(CARRYB_21__22_), .CI(SUMB_21__23_), .CO(
        CARRYB_22__22_), .S(SUMB_22__22_) );
  FA_X1 S2_22_23 ( .A(ab_22__23_), .B(CARRYB_21__23_), .CI(SUMB_21__24_), .CO(
        CARRYB_22__23_), .S(SUMB_22__23_) );
  FA_X1 S2_22_24 ( .A(ab_22__24_), .B(CARRYB_21__24_), .CI(SUMB_21__25_), .CO(
        CARRYB_22__24_), .S(SUMB_22__24_) );
  FA_X1 S2_22_25 ( .A(ab_22__25_), .B(CARRYB_21__25_), .CI(SUMB_21__26_), .CO(
        CARRYB_22__25_), .S(SUMB_22__25_) );
  FA_X1 S2_22_26 ( .A(ab_22__26_), .B(CARRYB_21__26_), .CI(SUMB_21__27_), .CO(
        CARRYB_22__26_), .S(SUMB_22__26_) );
  FA_X1 S2_22_27 ( .A(ab_22__27_), .B(CARRYB_21__27_), .CI(SUMB_21__28_), .CO(
        CARRYB_22__27_), .S(SUMB_22__27_) );
  FA_X1 S2_22_28 ( .A(ab_22__28_), .B(CARRYB_21__28_), .CI(SUMB_21__29_), .CO(
        CARRYB_22__28_), .S(SUMB_22__28_) );
  FA_X1 S2_22_29 ( .A(ab_22__29_), .B(CARRYB_21__29_), .CI(SUMB_21__30_), .CO(
        CARRYB_22__29_), .S(SUMB_22__29_) );
  FA_X1 S3_22_30 ( .A(ab_22__30_), .B(CARRYB_21__30_), .CI(ab_21__31_), .CO(
        CARRYB_22__30_), .S(SUMB_22__30_) );
  FA_X1 S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), .CO(
        CARRYB_21__0_), .S(A1_19_) );
  FA_X1 S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), .CO(
        CARRYB_21__1_), .S(SUMB_21__1_) );
  FA_X1 S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), .CO(
        CARRYB_21__2_), .S(SUMB_21__2_) );
  FA_X1 S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), .CO(
        CARRYB_21__3_), .S(SUMB_21__3_) );
  FA_X1 S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), .CO(
        CARRYB_21__4_), .S(SUMB_21__4_) );
  FA_X1 S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), .CO(
        CARRYB_21__5_), .S(SUMB_21__5_) );
  FA_X1 S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), .CO(
        CARRYB_21__6_), .S(SUMB_21__6_) );
  FA_X1 S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), .CO(
        CARRYB_21__7_), .S(SUMB_21__7_) );
  FA_X1 S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), .CO(
        CARRYB_21__8_), .S(SUMB_21__8_) );
  FA_X1 S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), .CO(
        CARRYB_21__9_), .S(SUMB_21__9_) );
  FA_X1 S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), .CO(
        CARRYB_21__10_), .S(SUMB_21__10_) );
  FA_X1 S2_21_11 ( .A(ab_21__11_), .B(CARRYB_20__11_), .CI(SUMB_20__12_), .CO(
        CARRYB_21__11_), .S(SUMB_21__11_) );
  FA_X1 S2_21_12 ( .A(ab_21__12_), .B(CARRYB_20__12_), .CI(SUMB_20__13_), .CO(
        CARRYB_21__12_), .S(SUMB_21__12_) );
  FA_X1 S2_21_13 ( .A(ab_21__13_), .B(CARRYB_20__13_), .CI(SUMB_20__14_), .CO(
        CARRYB_21__13_), .S(SUMB_21__13_) );
  FA_X1 S2_21_14 ( .A(ab_21__14_), .B(CARRYB_20__14_), .CI(SUMB_20__15_), .CO(
        CARRYB_21__14_), .S(SUMB_21__14_) );
  FA_X1 S2_21_15 ( .A(ab_21__15_), .B(CARRYB_20__15_), .CI(SUMB_20__16_), .CO(
        CARRYB_21__15_), .S(SUMB_21__15_) );
  FA_X1 S2_21_16 ( .A(ab_21__16_), .B(CARRYB_20__16_), .CI(SUMB_20__17_), .CO(
        CARRYB_21__16_), .S(SUMB_21__16_) );
  FA_X1 S2_21_17 ( .A(ab_21__17_), .B(CARRYB_20__17_), .CI(SUMB_20__18_), .CO(
        CARRYB_21__17_), .S(SUMB_21__17_) );
  FA_X1 S2_21_18 ( .A(ab_21__18_), .B(CARRYB_20__18_), .CI(SUMB_20__19_), .CO(
        CARRYB_21__18_), .S(SUMB_21__18_) );
  FA_X1 S2_21_19 ( .A(ab_21__19_), .B(CARRYB_20__19_), .CI(SUMB_20__20_), .CO(
        CARRYB_21__19_), .S(SUMB_21__19_) );
  FA_X1 S2_21_20 ( .A(ab_21__20_), .B(CARRYB_20__20_), .CI(SUMB_20__21_), .CO(
        CARRYB_21__20_), .S(SUMB_21__20_) );
  FA_X1 S2_21_21 ( .A(ab_21__21_), .B(CARRYB_20__21_), .CI(SUMB_20__22_), .CO(
        CARRYB_21__21_), .S(SUMB_21__21_) );
  FA_X1 S2_21_22 ( .A(ab_21__22_), .B(CARRYB_20__22_), .CI(SUMB_20__23_), .CO(
        CARRYB_21__22_), .S(SUMB_21__22_) );
  FA_X1 S2_21_23 ( .A(ab_21__23_), .B(CARRYB_20__23_), .CI(SUMB_20__24_), .CO(
        CARRYB_21__23_), .S(SUMB_21__23_) );
  FA_X1 S2_21_24 ( .A(ab_21__24_), .B(CARRYB_20__24_), .CI(SUMB_20__25_), .CO(
        CARRYB_21__24_), .S(SUMB_21__24_) );
  FA_X1 S2_21_25 ( .A(ab_21__25_), .B(CARRYB_20__25_), .CI(SUMB_20__26_), .CO(
        CARRYB_21__25_), .S(SUMB_21__25_) );
  FA_X1 S2_21_26 ( .A(ab_21__26_), .B(CARRYB_20__26_), .CI(SUMB_20__27_), .CO(
        CARRYB_21__26_), .S(SUMB_21__26_) );
  FA_X1 S2_21_27 ( .A(ab_21__27_), .B(CARRYB_20__27_), .CI(SUMB_20__28_), .CO(
        CARRYB_21__27_), .S(SUMB_21__27_) );
  FA_X1 S2_21_28 ( .A(ab_21__28_), .B(CARRYB_20__28_), .CI(SUMB_20__29_), .CO(
        CARRYB_21__28_), .S(SUMB_21__28_) );
  FA_X1 S2_21_29 ( .A(ab_21__29_), .B(CARRYB_20__29_), .CI(SUMB_20__30_), .CO(
        CARRYB_21__29_), .S(SUMB_21__29_) );
  FA_X1 S3_21_30 ( .A(ab_21__30_), .B(CARRYB_20__30_), .CI(ab_20__31_), .CO(
        CARRYB_21__30_), .S(SUMB_21__30_) );
  FA_X1 S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), .CO(
        CARRYB_20__0_), .S(A1_18_) );
  FA_X1 S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), .CO(
        CARRYB_20__1_), .S(SUMB_20__1_) );
  FA_X1 S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), .CO(
        CARRYB_20__2_), .S(SUMB_20__2_) );
  FA_X1 S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), .CO(
        CARRYB_20__3_), .S(SUMB_20__3_) );
  FA_X1 S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), .CO(
        CARRYB_20__4_), .S(SUMB_20__4_) );
  FA_X1 S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), .CO(
        CARRYB_20__5_), .S(SUMB_20__5_) );
  FA_X1 S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), .CO(
        CARRYB_20__6_), .S(SUMB_20__6_) );
  FA_X1 S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), .CO(
        CARRYB_20__7_), .S(SUMB_20__7_) );
  FA_X1 S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), .CO(
        CARRYB_20__8_), .S(SUMB_20__8_) );
  FA_X1 S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), .CO(
        CARRYB_20__9_), .S(SUMB_20__9_) );
  FA_X1 S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), .CO(
        CARRYB_20__10_), .S(SUMB_20__10_) );
  FA_X1 S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), .CO(
        CARRYB_20__11_), .S(SUMB_20__11_) );
  FA_X1 S2_20_12 ( .A(ab_20__12_), .B(CARRYB_19__12_), .CI(SUMB_19__13_), .CO(
        CARRYB_20__12_), .S(SUMB_20__12_) );
  FA_X1 S2_20_13 ( .A(ab_20__13_), .B(CARRYB_19__13_), .CI(SUMB_19__14_), .CO(
        CARRYB_20__13_), .S(SUMB_20__13_) );
  FA_X1 S2_20_14 ( .A(ab_20__14_), .B(CARRYB_19__14_), .CI(SUMB_19__15_), .CO(
        CARRYB_20__14_), .S(SUMB_20__14_) );
  FA_X1 S2_20_15 ( .A(ab_20__15_), .B(CARRYB_19__15_), .CI(SUMB_19__16_), .CO(
        CARRYB_20__15_), .S(SUMB_20__15_) );
  FA_X1 S2_20_16 ( .A(ab_20__16_), .B(CARRYB_19__16_), .CI(SUMB_19__17_), .CO(
        CARRYB_20__16_), .S(SUMB_20__16_) );
  FA_X1 S2_20_17 ( .A(ab_20__17_), .B(CARRYB_19__17_), .CI(SUMB_19__18_), .CO(
        CARRYB_20__17_), .S(SUMB_20__17_) );
  FA_X1 S2_20_18 ( .A(ab_20__18_), .B(CARRYB_19__18_), .CI(SUMB_19__19_), .CO(
        CARRYB_20__18_), .S(SUMB_20__18_) );
  FA_X1 S2_20_19 ( .A(ab_20__19_), .B(CARRYB_19__19_), .CI(SUMB_19__20_), .CO(
        CARRYB_20__19_), .S(SUMB_20__19_) );
  FA_X1 S2_20_20 ( .A(ab_20__20_), .B(CARRYB_19__20_), .CI(SUMB_19__21_), .CO(
        CARRYB_20__20_), .S(SUMB_20__20_) );
  FA_X1 S2_20_21 ( .A(ab_20__21_), .B(CARRYB_19__21_), .CI(SUMB_19__22_), .CO(
        CARRYB_20__21_), .S(SUMB_20__21_) );
  FA_X1 S2_20_22 ( .A(ab_20__22_), .B(CARRYB_19__22_), .CI(SUMB_19__23_), .CO(
        CARRYB_20__22_), .S(SUMB_20__22_) );
  FA_X1 S2_20_23 ( .A(ab_20__23_), .B(CARRYB_19__23_), .CI(SUMB_19__24_), .CO(
        CARRYB_20__23_), .S(SUMB_20__23_) );
  FA_X1 S2_20_24 ( .A(ab_20__24_), .B(CARRYB_19__24_), .CI(SUMB_19__25_), .CO(
        CARRYB_20__24_), .S(SUMB_20__24_) );
  FA_X1 S2_20_25 ( .A(ab_20__25_), .B(CARRYB_19__25_), .CI(SUMB_19__26_), .CO(
        CARRYB_20__25_), .S(SUMB_20__25_) );
  FA_X1 S2_20_26 ( .A(ab_20__26_), .B(CARRYB_19__26_), .CI(SUMB_19__27_), .CO(
        CARRYB_20__26_), .S(SUMB_20__26_) );
  FA_X1 S2_20_27 ( .A(ab_20__27_), .B(CARRYB_19__27_), .CI(SUMB_19__28_), .CO(
        CARRYB_20__27_), .S(SUMB_20__27_) );
  FA_X1 S2_20_28 ( .A(ab_20__28_), .B(CARRYB_19__28_), .CI(SUMB_19__29_), .CO(
        CARRYB_20__28_), .S(SUMB_20__28_) );
  FA_X1 S2_20_29 ( .A(ab_20__29_), .B(CARRYB_19__29_), .CI(SUMB_19__30_), .CO(
        CARRYB_20__29_), .S(SUMB_20__29_) );
  FA_X1 S3_20_30 ( .A(ab_20__30_), .B(CARRYB_19__30_), .CI(ab_19__31_), .CO(
        CARRYB_20__30_), .S(SUMB_20__30_) );
  FA_X1 S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), .CO(
        CARRYB_19__0_), .S(A1_17_) );
  FA_X1 S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), .CO(
        CARRYB_19__1_), .S(SUMB_19__1_) );
  FA_X1 S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), .CO(
        CARRYB_19__2_), .S(SUMB_19__2_) );
  FA_X1 S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), .CO(
        CARRYB_19__3_), .S(SUMB_19__3_) );
  FA_X1 S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), .CO(
        CARRYB_19__4_), .S(SUMB_19__4_) );
  FA_X1 S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), .CO(
        CARRYB_19__5_), .S(SUMB_19__5_) );
  FA_X1 S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), .CO(
        CARRYB_19__6_), .S(SUMB_19__6_) );
  FA_X1 S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), .CO(
        CARRYB_19__7_), .S(SUMB_19__7_) );
  FA_X1 S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), .CO(
        CARRYB_19__8_), .S(SUMB_19__8_) );
  FA_X1 S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), .CO(
        CARRYB_19__9_), .S(SUMB_19__9_) );
  FA_X1 S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), .CO(
        CARRYB_19__10_), .S(SUMB_19__10_) );
  FA_X1 S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), .CO(
        CARRYB_19__11_), .S(SUMB_19__11_) );
  FA_X1 S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), .CO(
        CARRYB_19__12_), .S(SUMB_19__12_) );
  FA_X1 S2_19_13 ( .A(ab_19__13_), .B(CARRYB_18__13_), .CI(SUMB_18__14_), .CO(
        CARRYB_19__13_), .S(SUMB_19__13_) );
  FA_X1 S2_19_14 ( .A(ab_19__14_), .B(CARRYB_18__14_), .CI(SUMB_18__15_), .CO(
        CARRYB_19__14_), .S(SUMB_19__14_) );
  FA_X1 S2_19_15 ( .A(ab_19__15_), .B(CARRYB_18__15_), .CI(SUMB_18__16_), .CO(
        CARRYB_19__15_), .S(SUMB_19__15_) );
  FA_X1 S2_19_16 ( .A(ab_19__16_), .B(CARRYB_18__16_), .CI(SUMB_18__17_), .CO(
        CARRYB_19__16_), .S(SUMB_19__16_) );
  FA_X1 S2_19_17 ( .A(ab_19__17_), .B(CARRYB_18__17_), .CI(SUMB_18__18_), .CO(
        CARRYB_19__17_), .S(SUMB_19__17_) );
  FA_X1 S2_19_18 ( .A(ab_19__18_), .B(CARRYB_18__18_), .CI(SUMB_18__19_), .CO(
        CARRYB_19__18_), .S(SUMB_19__18_) );
  FA_X1 S2_19_19 ( .A(ab_19__19_), .B(CARRYB_18__19_), .CI(SUMB_18__20_), .CO(
        CARRYB_19__19_), .S(SUMB_19__19_) );
  FA_X1 S2_19_20 ( .A(ab_19__20_), .B(CARRYB_18__20_), .CI(SUMB_18__21_), .CO(
        CARRYB_19__20_), .S(SUMB_19__20_) );
  FA_X1 S2_19_21 ( .A(ab_19__21_), .B(CARRYB_18__21_), .CI(SUMB_18__22_), .CO(
        CARRYB_19__21_), .S(SUMB_19__21_) );
  FA_X1 S2_19_22 ( .A(ab_19__22_), .B(CARRYB_18__22_), .CI(SUMB_18__23_), .CO(
        CARRYB_19__22_), .S(SUMB_19__22_) );
  FA_X1 S2_19_23 ( .A(ab_19__23_), .B(CARRYB_18__23_), .CI(SUMB_18__24_), .CO(
        CARRYB_19__23_), .S(SUMB_19__23_) );
  FA_X1 S2_19_24 ( .A(ab_19__24_), .B(CARRYB_18__24_), .CI(SUMB_18__25_), .CO(
        CARRYB_19__24_), .S(SUMB_19__24_) );
  FA_X1 S2_19_25 ( .A(ab_19__25_), .B(CARRYB_18__25_), .CI(SUMB_18__26_), .CO(
        CARRYB_19__25_), .S(SUMB_19__25_) );
  FA_X1 S2_19_26 ( .A(ab_19__26_), .B(CARRYB_18__26_), .CI(SUMB_18__27_), .CO(
        CARRYB_19__26_), .S(SUMB_19__26_) );
  FA_X1 S2_19_27 ( .A(ab_19__27_), .B(CARRYB_18__27_), .CI(SUMB_18__28_), .CO(
        CARRYB_19__27_), .S(SUMB_19__27_) );
  FA_X1 S2_19_28 ( .A(ab_19__28_), .B(CARRYB_18__28_), .CI(SUMB_18__29_), .CO(
        CARRYB_19__28_), .S(SUMB_19__28_) );
  FA_X1 S2_19_29 ( .A(ab_19__29_), .B(CARRYB_18__29_), .CI(SUMB_18__30_), .CO(
        CARRYB_19__29_), .S(SUMB_19__29_) );
  FA_X1 S3_19_30 ( .A(ab_19__30_), .B(CARRYB_18__30_), .CI(ab_18__31_), .CO(
        CARRYB_19__30_), .S(SUMB_19__30_) );
  FA_X1 S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), .CO(
        CARRYB_18__0_), .S(A1_16_) );
  FA_X1 S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), .CO(
        CARRYB_18__1_), .S(SUMB_18__1_) );
  FA_X1 S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), .CO(
        CARRYB_18__2_), .S(SUMB_18__2_) );
  FA_X1 S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), .CO(
        CARRYB_18__3_), .S(SUMB_18__3_) );
  FA_X1 S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), .CO(
        CARRYB_18__4_), .S(SUMB_18__4_) );
  FA_X1 S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), .CO(
        CARRYB_18__5_), .S(SUMB_18__5_) );
  FA_X1 S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), .CO(
        CARRYB_18__6_), .S(SUMB_18__6_) );
  FA_X1 S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), .CO(
        CARRYB_18__7_), .S(SUMB_18__7_) );
  FA_X1 S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), .CO(
        CARRYB_18__8_), .S(SUMB_18__8_) );
  FA_X1 S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), .CO(
        CARRYB_18__9_), .S(SUMB_18__9_) );
  FA_X1 S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), .CO(
        CARRYB_18__10_), .S(SUMB_18__10_) );
  FA_X1 S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), .CO(
        CARRYB_18__11_), .S(SUMB_18__11_) );
  FA_X1 S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), .CO(
        CARRYB_18__12_), .S(SUMB_18__12_) );
  FA_X1 S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), .CO(
        CARRYB_18__13_), .S(SUMB_18__13_) );
  FA_X1 S2_18_14 ( .A(ab_18__14_), .B(CARRYB_17__14_), .CI(SUMB_17__15_), .CO(
        CARRYB_18__14_), .S(SUMB_18__14_) );
  FA_X1 S2_18_15 ( .A(ab_18__15_), .B(CARRYB_17__15_), .CI(SUMB_17__16_), .CO(
        CARRYB_18__15_), .S(SUMB_18__15_) );
  FA_X1 S2_18_16 ( .A(ab_18__16_), .B(CARRYB_17__16_), .CI(SUMB_17__17_), .CO(
        CARRYB_18__16_), .S(SUMB_18__16_) );
  FA_X1 S2_18_17 ( .A(ab_18__17_), .B(CARRYB_17__17_), .CI(SUMB_17__18_), .CO(
        CARRYB_18__17_), .S(SUMB_18__17_) );
  FA_X1 S2_18_18 ( .A(ab_18__18_), .B(CARRYB_17__18_), .CI(SUMB_17__19_), .CO(
        CARRYB_18__18_), .S(SUMB_18__18_) );
  FA_X1 S2_18_19 ( .A(ab_18__19_), .B(CARRYB_17__19_), .CI(SUMB_17__20_), .CO(
        CARRYB_18__19_), .S(SUMB_18__19_) );
  FA_X1 S2_18_20 ( .A(ab_18__20_), .B(CARRYB_17__20_), .CI(SUMB_17__21_), .CO(
        CARRYB_18__20_), .S(SUMB_18__20_) );
  FA_X1 S2_18_21 ( .A(ab_18__21_), .B(CARRYB_17__21_), .CI(SUMB_17__22_), .CO(
        CARRYB_18__21_), .S(SUMB_18__21_) );
  FA_X1 S2_18_22 ( .A(ab_18__22_), .B(CARRYB_17__22_), .CI(SUMB_17__23_), .CO(
        CARRYB_18__22_), .S(SUMB_18__22_) );
  FA_X1 S2_18_23 ( .A(ab_18__23_), .B(CARRYB_17__23_), .CI(SUMB_17__24_), .CO(
        CARRYB_18__23_), .S(SUMB_18__23_) );
  FA_X1 S2_18_24 ( .A(ab_18__24_), .B(CARRYB_17__24_), .CI(SUMB_17__25_), .CO(
        CARRYB_18__24_), .S(SUMB_18__24_) );
  FA_X1 S2_18_25 ( .A(ab_18__25_), .B(CARRYB_17__25_), .CI(SUMB_17__26_), .CO(
        CARRYB_18__25_), .S(SUMB_18__25_) );
  FA_X1 S2_18_26 ( .A(ab_18__26_), .B(CARRYB_17__26_), .CI(SUMB_17__27_), .CO(
        CARRYB_18__26_), .S(SUMB_18__26_) );
  FA_X1 S2_18_27 ( .A(ab_18__27_), .B(CARRYB_17__27_), .CI(SUMB_17__28_), .CO(
        CARRYB_18__27_), .S(SUMB_18__27_) );
  FA_X1 S2_18_28 ( .A(ab_18__28_), .B(CARRYB_17__28_), .CI(SUMB_17__29_), .CO(
        CARRYB_18__28_), .S(SUMB_18__28_) );
  FA_X1 S2_18_29 ( .A(ab_18__29_), .B(CARRYB_17__29_), .CI(SUMB_17__30_), .CO(
        CARRYB_18__29_), .S(SUMB_18__29_) );
  FA_X1 S3_18_30 ( .A(ab_18__30_), .B(CARRYB_17__30_), .CI(ab_17__31_), .CO(
        CARRYB_18__30_), .S(SUMB_18__30_) );
  FA_X1 S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), .CO(
        CARRYB_17__0_), .S(A1_15_) );
  FA_X1 S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), .CO(
        CARRYB_17__1_), .S(SUMB_17__1_) );
  FA_X1 S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), .CO(
        CARRYB_17__2_), .S(SUMB_17__2_) );
  FA_X1 S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), .CO(
        CARRYB_17__3_), .S(SUMB_17__3_) );
  FA_X1 S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), .CO(
        CARRYB_17__4_), .S(SUMB_17__4_) );
  FA_X1 S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), .CO(
        CARRYB_17__5_), .S(SUMB_17__5_) );
  FA_X1 S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), .CO(
        CARRYB_17__6_), .S(SUMB_17__6_) );
  FA_X1 S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), .CO(
        CARRYB_17__7_), .S(SUMB_17__7_) );
  FA_X1 S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), .CO(
        CARRYB_17__8_), .S(SUMB_17__8_) );
  FA_X1 S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), .CO(
        CARRYB_17__9_), .S(SUMB_17__9_) );
  FA_X1 S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), .CO(
        CARRYB_17__10_), .S(SUMB_17__10_) );
  FA_X1 S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), .CO(
        CARRYB_17__11_), .S(SUMB_17__11_) );
  FA_X1 S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), .CO(
        CARRYB_17__12_), .S(SUMB_17__12_) );
  FA_X1 S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), .CO(
        CARRYB_17__13_), .S(SUMB_17__13_) );
  FA_X1 S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), .CO(
        CARRYB_17__14_), .S(SUMB_17__14_) );
  FA_X1 S2_17_15 ( .A(ab_17__15_), .B(CARRYB_16__15_), .CI(SUMB_16__16_), .CO(
        CARRYB_17__15_), .S(SUMB_17__15_) );
  FA_X1 S2_17_16 ( .A(ab_17__16_), .B(CARRYB_16__16_), .CI(SUMB_16__17_), .CO(
        CARRYB_17__16_), .S(SUMB_17__16_) );
  FA_X1 S2_17_17 ( .A(ab_17__17_), .B(CARRYB_16__17_), .CI(SUMB_16__18_), .CO(
        CARRYB_17__17_), .S(SUMB_17__17_) );
  FA_X1 S2_17_18 ( .A(ab_17__18_), .B(CARRYB_16__18_), .CI(SUMB_16__19_), .CO(
        CARRYB_17__18_), .S(SUMB_17__18_) );
  FA_X1 S2_17_19 ( .A(ab_17__19_), .B(CARRYB_16__19_), .CI(SUMB_16__20_), .CO(
        CARRYB_17__19_), .S(SUMB_17__19_) );
  FA_X1 S2_17_20 ( .A(ab_17__20_), .B(CARRYB_16__20_), .CI(SUMB_16__21_), .CO(
        CARRYB_17__20_), .S(SUMB_17__20_) );
  FA_X1 S2_17_21 ( .A(ab_17__21_), .B(CARRYB_16__21_), .CI(SUMB_16__22_), .CO(
        CARRYB_17__21_), .S(SUMB_17__21_) );
  FA_X1 S2_17_22 ( .A(ab_17__22_), .B(CARRYB_16__22_), .CI(SUMB_16__23_), .CO(
        CARRYB_17__22_), .S(SUMB_17__22_) );
  FA_X1 S2_17_23 ( .A(ab_17__23_), .B(CARRYB_16__23_), .CI(SUMB_16__24_), .CO(
        CARRYB_17__23_), .S(SUMB_17__23_) );
  FA_X1 S2_17_24 ( .A(ab_17__24_), .B(CARRYB_16__24_), .CI(SUMB_16__25_), .CO(
        CARRYB_17__24_), .S(SUMB_17__24_) );
  FA_X1 S2_17_25 ( .A(ab_17__25_), .B(CARRYB_16__25_), .CI(SUMB_16__26_), .CO(
        CARRYB_17__25_), .S(SUMB_17__25_) );
  FA_X1 S2_17_26 ( .A(ab_17__26_), .B(CARRYB_16__26_), .CI(SUMB_16__27_), .CO(
        CARRYB_17__26_), .S(SUMB_17__26_) );
  FA_X1 S2_17_27 ( .A(ab_17__27_), .B(CARRYB_16__27_), .CI(SUMB_16__28_), .CO(
        CARRYB_17__27_), .S(SUMB_17__27_) );
  FA_X1 S2_17_28 ( .A(ab_17__28_), .B(CARRYB_16__28_), .CI(SUMB_16__29_), .CO(
        CARRYB_17__28_), .S(SUMB_17__28_) );
  FA_X1 S2_17_29 ( .A(ab_17__29_), .B(CARRYB_16__29_), .CI(SUMB_16__30_), .CO(
        CARRYB_17__29_), .S(SUMB_17__29_) );
  FA_X1 S3_17_30 ( .A(ab_17__30_), .B(CARRYB_16__30_), .CI(ab_16__31_), .CO(
        CARRYB_17__30_), .S(SUMB_17__30_) );
  FA_X1 S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(A1_14_) );
  FA_X1 S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  FA_X1 S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  FA_X1 S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  FA_X1 S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  FA_X1 S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  FA_X1 S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  FA_X1 S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), .CO(
        CARRYB_16__7_), .S(SUMB_16__7_) );
  FA_X1 S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), .CO(
        CARRYB_16__8_), .S(SUMB_16__8_) );
  FA_X1 S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), .CO(
        CARRYB_16__9_), .S(SUMB_16__9_) );
  FA_X1 S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), .CO(
        CARRYB_16__10_), .S(SUMB_16__10_) );
  FA_X1 S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), .CO(
        CARRYB_16__11_), .S(SUMB_16__11_) );
  FA_X1 S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), .CO(
        CARRYB_16__12_), .S(SUMB_16__12_) );
  FA_X1 S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), .CO(
        CARRYB_16__13_), .S(SUMB_16__13_) );
  FA_X1 S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), .CO(
        CARRYB_16__14_), .S(SUMB_16__14_) );
  FA_X1 S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), .CO(
        CARRYB_16__15_), .S(SUMB_16__15_) );
  FA_X1 S2_16_16 ( .A(ab_16__16_), .B(CARRYB_15__16_), .CI(SUMB_15__17_), .CO(
        CARRYB_16__16_), .S(SUMB_16__16_) );
  FA_X1 S2_16_17 ( .A(ab_16__17_), .B(CARRYB_15__17_), .CI(SUMB_15__18_), .CO(
        CARRYB_16__17_), .S(SUMB_16__17_) );
  FA_X1 S2_16_18 ( .A(ab_16__18_), .B(CARRYB_15__18_), .CI(SUMB_15__19_), .CO(
        CARRYB_16__18_), .S(SUMB_16__18_) );
  FA_X1 S2_16_19 ( .A(ab_16__19_), .B(CARRYB_15__19_), .CI(SUMB_15__20_), .CO(
        CARRYB_16__19_), .S(SUMB_16__19_) );
  FA_X1 S2_16_20 ( .A(ab_16__20_), .B(CARRYB_15__20_), .CI(SUMB_15__21_), .CO(
        CARRYB_16__20_), .S(SUMB_16__20_) );
  FA_X1 S2_16_21 ( .A(ab_16__21_), .B(CARRYB_15__21_), .CI(SUMB_15__22_), .CO(
        CARRYB_16__21_), .S(SUMB_16__21_) );
  FA_X1 S2_16_22 ( .A(ab_16__22_), .B(CARRYB_15__22_), .CI(SUMB_15__23_), .CO(
        CARRYB_16__22_), .S(SUMB_16__22_) );
  FA_X1 S2_16_23 ( .A(ab_16__23_), .B(CARRYB_15__23_), .CI(SUMB_15__24_), .CO(
        CARRYB_16__23_), .S(SUMB_16__23_) );
  FA_X1 S2_16_24 ( .A(ab_16__24_), .B(CARRYB_15__24_), .CI(SUMB_15__25_), .CO(
        CARRYB_16__24_), .S(SUMB_16__24_) );
  FA_X1 S2_16_25 ( .A(ab_16__25_), .B(CARRYB_15__25_), .CI(SUMB_15__26_), .CO(
        CARRYB_16__25_), .S(SUMB_16__25_) );
  FA_X1 S2_16_26 ( .A(ab_16__26_), .B(CARRYB_15__26_), .CI(SUMB_15__27_), .CO(
        CARRYB_16__26_), .S(SUMB_16__26_) );
  FA_X1 S2_16_27 ( .A(ab_16__27_), .B(CARRYB_15__27_), .CI(SUMB_15__28_), .CO(
        CARRYB_16__27_), .S(SUMB_16__27_) );
  FA_X1 S2_16_28 ( .A(ab_16__28_), .B(CARRYB_15__28_), .CI(SUMB_15__29_), .CO(
        CARRYB_16__28_), .S(SUMB_16__28_) );
  FA_X1 S2_16_29 ( .A(ab_16__29_), .B(CARRYB_15__29_), .CI(SUMB_15__30_), .CO(
        CARRYB_16__29_), .S(SUMB_16__29_) );
  FA_X1 S3_16_30 ( .A(ab_16__30_), .B(CARRYB_15__30_), .CI(ab_15__31_), .CO(
        CARRYB_16__30_), .S(SUMB_16__30_) );
  FA_X1 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  FA_X1 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  FA_X1 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  FA_X1 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  FA_X1 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  FA_X1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  FA_X1 S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  FA_X1 S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  FA_X1 S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  FA_X1 S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  FA_X1 S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), .CO(
        CARRYB_15__10_), .S(SUMB_15__10_) );
  FA_X1 S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), .CO(
        CARRYB_15__11_), .S(SUMB_15__11_) );
  FA_X1 S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), .CO(
        CARRYB_15__12_), .S(SUMB_15__12_) );
  FA_X1 S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), .CO(
        CARRYB_15__13_), .S(SUMB_15__13_) );
  FA_X1 S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), .CO(
        CARRYB_15__14_), .S(SUMB_15__14_) );
  FA_X1 S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  FA_X1 S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), .CO(
        CARRYB_15__16_), .S(SUMB_15__16_) );
  FA_X1 S2_15_17 ( .A(ab_15__17_), .B(CARRYB_14__17_), .CI(SUMB_14__18_), .CO(
        CARRYB_15__17_), .S(SUMB_15__17_) );
  FA_X1 S2_15_18 ( .A(ab_15__18_), .B(CARRYB_14__18_), .CI(SUMB_14__19_), .CO(
        CARRYB_15__18_), .S(SUMB_15__18_) );
  FA_X1 S2_15_19 ( .A(ab_15__19_), .B(CARRYB_14__19_), .CI(SUMB_14__20_), .CO(
        CARRYB_15__19_), .S(SUMB_15__19_) );
  FA_X1 S2_15_20 ( .A(ab_15__20_), .B(CARRYB_14__20_), .CI(SUMB_14__21_), .CO(
        CARRYB_15__20_), .S(SUMB_15__20_) );
  FA_X1 S2_15_21 ( .A(ab_15__21_), .B(CARRYB_14__21_), .CI(SUMB_14__22_), .CO(
        CARRYB_15__21_), .S(SUMB_15__21_) );
  FA_X1 S2_15_22 ( .A(ab_15__22_), .B(CARRYB_14__22_), .CI(SUMB_14__23_), .CO(
        CARRYB_15__22_), .S(SUMB_15__22_) );
  FA_X1 S2_15_23 ( .A(ab_15__23_), .B(CARRYB_14__23_), .CI(SUMB_14__24_), .CO(
        CARRYB_15__23_), .S(SUMB_15__23_) );
  FA_X1 S2_15_24 ( .A(ab_15__24_), .B(CARRYB_14__24_), .CI(SUMB_14__25_), .CO(
        CARRYB_15__24_), .S(SUMB_15__24_) );
  FA_X1 S2_15_25 ( .A(ab_15__25_), .B(CARRYB_14__25_), .CI(SUMB_14__26_), .CO(
        CARRYB_15__25_), .S(SUMB_15__25_) );
  FA_X1 S2_15_26 ( .A(ab_15__26_), .B(CARRYB_14__26_), .CI(SUMB_14__27_), .CO(
        CARRYB_15__26_), .S(SUMB_15__26_) );
  FA_X1 S2_15_27 ( .A(ab_15__27_), .B(CARRYB_14__27_), .CI(SUMB_14__28_), .CO(
        CARRYB_15__27_), .S(SUMB_15__27_) );
  FA_X1 S2_15_28 ( .A(ab_15__28_), .B(CARRYB_14__28_), .CI(SUMB_14__29_), .CO(
        CARRYB_15__28_), .S(SUMB_15__28_) );
  FA_X1 S2_15_29 ( .A(ab_15__29_), .B(CARRYB_14__29_), .CI(SUMB_14__30_), .CO(
        CARRYB_15__29_), .S(SUMB_15__29_) );
  FA_X1 S3_15_30 ( .A(ab_15__30_), .B(CARRYB_14__30_), .CI(ab_14__31_), .CO(
        CARRYB_15__30_), .S(SUMB_15__30_) );
  FA_X1 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  FA_X1 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  FA_X1 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  FA_X1 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  FA_X1 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  FA_X1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  FA_X1 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  FA_X1 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  FA_X1 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  FA_X1 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  FA_X1 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), .CO(
        CARRYB_14__10_), .S(SUMB_14__10_) );
  FA_X1 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), .CO(
        CARRYB_14__11_), .S(SUMB_14__11_) );
  FA_X1 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), .CO(
        CARRYB_14__12_), .S(SUMB_14__12_) );
  FA_X1 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), .CO(
        CARRYB_14__13_), .S(SUMB_14__13_) );
  FA_X1 S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  FA_X1 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), .CO(
        CARRYB_14__15_), .S(SUMB_14__15_) );
  FA_X1 S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), .CO(
        CARRYB_14__16_), .S(SUMB_14__16_) );
  FA_X1 S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), .CO(
        CARRYB_14__17_), .S(SUMB_14__17_) );
  FA_X1 S2_14_18 ( .A(ab_14__18_), .B(CARRYB_13__18_), .CI(SUMB_13__19_), .CO(
        CARRYB_14__18_), .S(SUMB_14__18_) );
  FA_X1 S2_14_19 ( .A(ab_14__19_), .B(CARRYB_13__19_), .CI(SUMB_13__20_), .CO(
        CARRYB_14__19_), .S(SUMB_14__19_) );
  FA_X1 S2_14_20 ( .A(ab_14__20_), .B(CARRYB_13__20_), .CI(SUMB_13__21_), .CO(
        CARRYB_14__20_), .S(SUMB_14__20_) );
  FA_X1 S2_14_21 ( .A(ab_14__21_), .B(CARRYB_13__21_), .CI(SUMB_13__22_), .CO(
        CARRYB_14__21_), .S(SUMB_14__21_) );
  FA_X1 S2_14_22 ( .A(ab_14__22_), .B(CARRYB_13__22_), .CI(SUMB_13__23_), .CO(
        CARRYB_14__22_), .S(SUMB_14__22_) );
  FA_X1 S2_14_23 ( .A(ab_14__23_), .B(CARRYB_13__23_), .CI(SUMB_13__24_), .CO(
        CARRYB_14__23_), .S(SUMB_14__23_) );
  FA_X1 S2_14_24 ( .A(ab_14__24_), .B(CARRYB_13__24_), .CI(SUMB_13__25_), .CO(
        CARRYB_14__24_), .S(SUMB_14__24_) );
  FA_X1 S2_14_25 ( .A(ab_14__25_), .B(CARRYB_13__25_), .CI(SUMB_13__26_), .CO(
        CARRYB_14__25_), .S(SUMB_14__25_) );
  FA_X1 S2_14_26 ( .A(ab_14__26_), .B(CARRYB_13__26_), .CI(SUMB_13__27_), .CO(
        CARRYB_14__26_), .S(SUMB_14__26_) );
  FA_X1 S2_14_27 ( .A(ab_14__27_), .B(CARRYB_13__27_), .CI(SUMB_13__28_), .CO(
        CARRYB_14__27_), .S(SUMB_14__27_) );
  FA_X1 S2_14_28 ( .A(ab_14__28_), .B(CARRYB_13__28_), .CI(SUMB_13__29_), .CO(
        CARRYB_14__28_), .S(SUMB_14__28_) );
  FA_X1 S2_14_29 ( .A(ab_14__29_), .B(CARRYB_13__29_), .CI(SUMB_13__30_), .CO(
        CARRYB_14__29_), .S(SUMB_14__29_) );
  FA_X1 S3_14_30 ( .A(ab_14__30_), .B(CARRYB_13__30_), .CI(ab_13__31_), .CO(
        CARRYB_14__30_), .S(SUMB_14__30_) );
  FA_X1 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  FA_X1 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  FA_X1 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  FA_X1 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  FA_X1 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  FA_X1 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  FA_X1 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  FA_X1 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  FA_X1 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  FA_X1 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  FA_X1 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), .CO(
        CARRYB_13__10_), .S(SUMB_13__10_) );
  FA_X1 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), .CO(
        CARRYB_13__11_), .S(SUMB_13__11_) );
  FA_X1 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), .CO(
        CARRYB_13__12_), .S(SUMB_13__12_) );
  FA_X1 S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  FA_X1 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), .CO(
        CARRYB_13__14_), .S(SUMB_13__14_) );
  FA_X1 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), .CO(
        CARRYB_13__15_), .S(SUMB_13__15_) );
  FA_X1 S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), .CO(
        CARRYB_13__16_), .S(SUMB_13__16_) );
  FA_X1 S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), .CO(
        CARRYB_13__17_), .S(SUMB_13__17_) );
  FA_X1 S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), .CO(
        CARRYB_13__18_), .S(SUMB_13__18_) );
  FA_X1 S2_13_19 ( .A(ab_13__19_), .B(CARRYB_12__19_), .CI(SUMB_12__20_), .CO(
        CARRYB_13__19_), .S(SUMB_13__19_) );
  FA_X1 S2_13_20 ( .A(ab_13__20_), .B(CARRYB_12__20_), .CI(SUMB_12__21_), .CO(
        CARRYB_13__20_), .S(SUMB_13__20_) );
  FA_X1 S2_13_21 ( .A(ab_13__21_), .B(CARRYB_12__21_), .CI(SUMB_12__22_), .CO(
        CARRYB_13__21_), .S(SUMB_13__21_) );
  FA_X1 S2_13_22 ( .A(ab_13__22_), .B(CARRYB_12__22_), .CI(SUMB_12__23_), .CO(
        CARRYB_13__22_), .S(SUMB_13__22_) );
  FA_X1 S2_13_23 ( .A(ab_13__23_), .B(CARRYB_12__23_), .CI(SUMB_12__24_), .CO(
        CARRYB_13__23_), .S(SUMB_13__23_) );
  FA_X1 S2_13_24 ( .A(ab_13__24_), .B(CARRYB_12__24_), .CI(SUMB_12__25_), .CO(
        CARRYB_13__24_), .S(SUMB_13__24_) );
  FA_X1 S2_13_25 ( .A(ab_13__25_), .B(CARRYB_12__25_), .CI(SUMB_12__26_), .CO(
        CARRYB_13__25_), .S(SUMB_13__25_) );
  FA_X1 S2_13_26 ( .A(ab_13__26_), .B(CARRYB_12__26_), .CI(SUMB_12__27_), .CO(
        CARRYB_13__26_), .S(SUMB_13__26_) );
  FA_X1 S2_13_27 ( .A(ab_13__27_), .B(CARRYB_12__27_), .CI(SUMB_12__28_), .CO(
        CARRYB_13__27_), .S(SUMB_13__27_) );
  FA_X1 S2_13_28 ( .A(ab_13__28_), .B(CARRYB_12__28_), .CI(SUMB_12__29_), .CO(
        CARRYB_13__28_), .S(SUMB_13__28_) );
  FA_X1 S2_13_29 ( .A(ab_13__29_), .B(CARRYB_12__29_), .CI(SUMB_12__30_), .CO(
        CARRYB_13__29_), .S(SUMB_13__29_) );
  FA_X1 S3_13_30 ( .A(ab_13__30_), .B(CARRYB_12__30_), .CI(ab_12__31_), .CO(
        CARRYB_13__30_), .S(SUMB_13__30_) );
  FA_X1 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  FA_X1 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  FA_X1 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  FA_X1 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  FA_X1 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  FA_X1 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  FA_X1 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  FA_X1 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  FA_X1 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  FA_X1 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  FA_X1 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), .CO(
        CARRYB_12__10_), .S(SUMB_12__10_) );
  FA_X1 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), .CO(
        CARRYB_12__11_), .S(SUMB_12__11_) );
  FA_X1 S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  FA_X1 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), .CO(
        CARRYB_12__13_), .S(SUMB_12__13_) );
  FA_X1 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), .CO(
        CARRYB_12__14_), .S(SUMB_12__14_) );
  FA_X1 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), .CO(
        CARRYB_12__15_), .S(SUMB_12__15_) );
  FA_X1 S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), .CO(
        CARRYB_12__16_), .S(SUMB_12__16_) );
  FA_X1 S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), .CO(
        CARRYB_12__17_), .S(SUMB_12__17_) );
  FA_X1 S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), .CO(
        CARRYB_12__18_), .S(SUMB_12__18_) );
  FA_X1 S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), .CO(
        CARRYB_12__19_), .S(SUMB_12__19_) );
  FA_X1 S2_12_20 ( .A(ab_12__20_), .B(CARRYB_11__20_), .CI(SUMB_11__21_), .CO(
        CARRYB_12__20_), .S(SUMB_12__20_) );
  FA_X1 S2_12_21 ( .A(ab_12__21_), .B(CARRYB_11__21_), .CI(SUMB_11__22_), .CO(
        CARRYB_12__21_), .S(SUMB_12__21_) );
  FA_X1 S2_12_22 ( .A(ab_12__22_), .B(CARRYB_11__22_), .CI(SUMB_11__23_), .CO(
        CARRYB_12__22_), .S(SUMB_12__22_) );
  FA_X1 S2_12_23 ( .A(ab_12__23_), .B(CARRYB_11__23_), .CI(SUMB_11__24_), .CO(
        CARRYB_12__23_), .S(SUMB_12__23_) );
  FA_X1 S2_12_24 ( .A(ab_12__24_), .B(CARRYB_11__24_), .CI(SUMB_11__25_), .CO(
        CARRYB_12__24_), .S(SUMB_12__24_) );
  FA_X1 S2_12_25 ( .A(ab_12__25_), .B(CARRYB_11__25_), .CI(SUMB_11__26_), .CO(
        CARRYB_12__25_), .S(SUMB_12__25_) );
  FA_X1 S2_12_26 ( .A(ab_12__26_), .B(CARRYB_11__26_), .CI(SUMB_11__27_), .CO(
        CARRYB_12__26_), .S(SUMB_12__26_) );
  FA_X1 S2_12_27 ( .A(ab_12__27_), .B(CARRYB_11__27_), .CI(SUMB_11__28_), .CO(
        CARRYB_12__27_), .S(SUMB_12__27_) );
  FA_X1 S2_12_28 ( .A(ab_12__28_), .B(CARRYB_11__28_), .CI(SUMB_11__29_), .CO(
        CARRYB_12__28_), .S(SUMB_12__28_) );
  FA_X1 S2_12_29 ( .A(ab_12__29_), .B(CARRYB_11__29_), .CI(SUMB_11__30_), .CO(
        CARRYB_12__29_), .S(SUMB_12__29_) );
  FA_X1 S3_12_30 ( .A(ab_12__30_), .B(CARRYB_11__30_), .CI(ab_11__31_), .CO(
        CARRYB_12__30_), .S(SUMB_12__30_) );
  FA_X1 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  FA_X1 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  FA_X1 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  FA_X1 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  FA_X1 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  FA_X1 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  FA_X1 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  FA_X1 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  FA_X1 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  FA_X1 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  FA_X1 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), .CO(
        CARRYB_11__10_), .S(SUMB_11__10_) );
  FA_X1 S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  FA_X1 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), .CO(
        CARRYB_11__12_), .S(SUMB_11__12_) );
  FA_X1 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), .CO(
        CARRYB_11__13_), .S(SUMB_11__13_) );
  FA_X1 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), .CO(
        CARRYB_11__14_), .S(SUMB_11__14_) );
  FA_X1 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), .CO(
        CARRYB_11__15_), .S(SUMB_11__15_) );
  FA_X1 S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), .CO(
        CARRYB_11__16_), .S(SUMB_11__16_) );
  FA_X1 S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), .CO(
        CARRYB_11__17_), .S(SUMB_11__17_) );
  FA_X1 S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), .CO(
        CARRYB_11__18_), .S(SUMB_11__18_) );
  FA_X1 S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), .CO(
        CARRYB_11__19_), .S(SUMB_11__19_) );
  FA_X1 S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), .CO(
        CARRYB_11__20_), .S(SUMB_11__20_) );
  FA_X1 S2_11_21 ( .A(ab_11__21_), .B(CARRYB_10__21_), .CI(SUMB_10__22_), .CO(
        CARRYB_11__21_), .S(SUMB_11__21_) );
  FA_X1 S2_11_22 ( .A(ab_11__22_), .B(CARRYB_10__22_), .CI(SUMB_10__23_), .CO(
        CARRYB_11__22_), .S(SUMB_11__22_) );
  FA_X1 S2_11_23 ( .A(ab_11__23_), .B(CARRYB_10__23_), .CI(SUMB_10__24_), .CO(
        CARRYB_11__23_), .S(SUMB_11__23_) );
  FA_X1 S2_11_24 ( .A(ab_11__24_), .B(CARRYB_10__24_), .CI(SUMB_10__25_), .CO(
        CARRYB_11__24_), .S(SUMB_11__24_) );
  FA_X1 S2_11_25 ( .A(ab_11__25_), .B(CARRYB_10__25_), .CI(SUMB_10__26_), .CO(
        CARRYB_11__25_), .S(SUMB_11__25_) );
  FA_X1 S2_11_26 ( .A(ab_11__26_), .B(CARRYB_10__26_), .CI(SUMB_10__27_), .CO(
        CARRYB_11__26_), .S(SUMB_11__26_) );
  FA_X1 S2_11_27 ( .A(ab_11__27_), .B(CARRYB_10__27_), .CI(SUMB_10__28_), .CO(
        CARRYB_11__27_), .S(SUMB_11__27_) );
  FA_X1 S2_11_28 ( .A(ab_11__28_), .B(CARRYB_10__28_), .CI(SUMB_10__29_), .CO(
        CARRYB_11__28_), .S(SUMB_11__28_) );
  FA_X1 S2_11_29 ( .A(ab_11__29_), .B(CARRYB_10__29_), .CI(SUMB_10__30_), .CO(
        CARRYB_11__29_), .S(SUMB_11__29_) );
  FA_X1 S3_11_30 ( .A(ab_11__30_), .B(CARRYB_10__30_), .CI(ab_10__31_), .CO(
        CARRYB_11__30_), .S(SUMB_11__30_) );
  FA_X1 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  FA_X1 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FA_X1 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FA_X1 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FA_X1 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FA_X1 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FA_X1 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FA_X1 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FA_X1 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FA_X1 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FA_X1 S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  FA_X1 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  FA_X1 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  FA_X1 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  FA_X1 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  FA_X1 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  FA_X1 S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  FA_X1 S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), .CO(
        CARRYB_10__17_), .S(SUMB_10__17_) );
  FA_X1 S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), .CO(
        CARRYB_10__18_), .S(SUMB_10__18_) );
  FA_X1 S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), .CO(
        CARRYB_10__19_), .S(SUMB_10__19_) );
  FA_X1 S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), .CO(
        CARRYB_10__20_), .S(SUMB_10__20_) );
  FA_X1 S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), .CO(
        CARRYB_10__21_), .S(SUMB_10__21_) );
  FA_X1 S2_10_22 ( .A(ab_10__22_), .B(CARRYB_9__22_), .CI(SUMB_9__23_), .CO(
        CARRYB_10__22_), .S(SUMB_10__22_) );
  FA_X1 S2_10_23 ( .A(ab_10__23_), .B(CARRYB_9__23_), .CI(SUMB_9__24_), .CO(
        CARRYB_10__23_), .S(SUMB_10__23_) );
  FA_X1 S2_10_24 ( .A(ab_10__24_), .B(CARRYB_9__24_), .CI(SUMB_9__25_), .CO(
        CARRYB_10__24_), .S(SUMB_10__24_) );
  FA_X1 S2_10_25 ( .A(ab_10__25_), .B(CARRYB_9__25_), .CI(SUMB_9__26_), .CO(
        CARRYB_10__25_), .S(SUMB_10__25_) );
  FA_X1 S2_10_26 ( .A(ab_10__26_), .B(CARRYB_9__26_), .CI(SUMB_9__27_), .CO(
        CARRYB_10__26_), .S(SUMB_10__26_) );
  FA_X1 S2_10_27 ( .A(ab_10__27_), .B(CARRYB_9__27_), .CI(SUMB_9__28_), .CO(
        CARRYB_10__27_), .S(SUMB_10__27_) );
  FA_X1 S2_10_28 ( .A(ab_10__28_), .B(CARRYB_9__28_), .CI(SUMB_9__29_), .CO(
        CARRYB_10__28_), .S(SUMB_10__28_) );
  FA_X1 S2_10_29 ( .A(ab_10__29_), .B(CARRYB_9__29_), .CI(SUMB_9__30_), .CO(
        CARRYB_10__29_), .S(SUMB_10__29_) );
  FA_X1 S3_10_30 ( .A(ab_10__30_), .B(CARRYB_9__30_), .CI(ab_9__31_), .CO(
        CARRYB_10__30_), .S(SUMB_10__30_) );
  FA_X1 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  FA_X1 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FA_X1 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FA_X1 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FA_X1 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FA_X1 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FA_X1 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FA_X1 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FA_X1 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FA_X1 S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FA_X1 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  FA_X1 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  FA_X1 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  FA_X1 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  FA_X1 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  FA_X1 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  FA_X1 S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  FA_X1 S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), .CO(
        CARRYB_9__17_), .S(SUMB_9__17_) );
  FA_X1 S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), .CO(
        CARRYB_9__18_), .S(SUMB_9__18_) );
  FA_X1 S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), .CO(
        CARRYB_9__19_), .S(SUMB_9__19_) );
  FA_X1 S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), .CO(
        CARRYB_9__20_), .S(SUMB_9__20_) );
  FA_X1 S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), .CO(
        CARRYB_9__21_), .S(SUMB_9__21_) );
  FA_X1 S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(SUMB_8__23_), .CO(
        CARRYB_9__22_), .S(SUMB_9__22_) );
  FA_X1 S2_9_23 ( .A(ab_9__23_), .B(CARRYB_8__23_), .CI(SUMB_8__24_), .CO(
        CARRYB_9__23_), .S(SUMB_9__23_) );
  FA_X1 S2_9_24 ( .A(ab_9__24_), .B(CARRYB_8__24_), .CI(SUMB_8__25_), .CO(
        CARRYB_9__24_), .S(SUMB_9__24_) );
  FA_X1 S2_9_25 ( .A(ab_9__25_), .B(CARRYB_8__25_), .CI(SUMB_8__26_), .CO(
        CARRYB_9__25_), .S(SUMB_9__25_) );
  FA_X1 S2_9_26 ( .A(ab_9__26_), .B(CARRYB_8__26_), .CI(SUMB_8__27_), .CO(
        CARRYB_9__26_), .S(SUMB_9__26_) );
  FA_X1 S2_9_27 ( .A(ab_9__27_), .B(CARRYB_8__27_), .CI(SUMB_8__28_), .CO(
        CARRYB_9__27_), .S(SUMB_9__27_) );
  FA_X1 S2_9_28 ( .A(ab_9__28_), .B(CARRYB_8__28_), .CI(SUMB_8__29_), .CO(
        CARRYB_9__28_), .S(SUMB_9__28_) );
  FA_X1 S2_9_29 ( .A(ab_9__29_), .B(CARRYB_8__29_), .CI(SUMB_8__30_), .CO(
        CARRYB_9__29_), .S(SUMB_9__29_) );
  FA_X1 S3_9_30 ( .A(ab_9__30_), .B(CARRYB_8__30_), .CI(ab_8__31_), .CO(
        CARRYB_9__30_), .S(SUMB_9__30_) );
  FA_X1 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  FA_X1 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FA_X1 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FA_X1 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FA_X1 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FA_X1 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FA_X1 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FA_X1 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FA_X1 S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FA_X1 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FA_X1 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  FA_X1 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  FA_X1 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  FA_X1 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  FA_X1 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  FA_X1 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  FA_X1 S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  FA_X1 S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), .CO(
        CARRYB_8__17_), .S(SUMB_8__17_) );
  FA_X1 S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), .CO(
        CARRYB_8__18_), .S(SUMB_8__18_) );
  FA_X1 S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), .CO(
        CARRYB_8__19_), .S(SUMB_8__19_) );
  FA_X1 S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), .CO(
        CARRYB_8__20_), .S(SUMB_8__20_) );
  FA_X1 S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), .CO(
        CARRYB_8__21_), .S(SUMB_8__21_) );
  FA_X1 S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), .CO(
        CARRYB_8__22_), .S(SUMB_8__22_) );
  FA_X1 S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .CI(SUMB_7__24_), .CO(
        CARRYB_8__23_), .S(SUMB_8__23_) );
  FA_X1 S2_8_24 ( .A(ab_8__24_), .B(CARRYB_7__24_), .CI(SUMB_7__25_), .CO(
        CARRYB_8__24_), .S(SUMB_8__24_) );
  FA_X1 S2_8_25 ( .A(ab_8__25_), .B(CARRYB_7__25_), .CI(SUMB_7__26_), .CO(
        CARRYB_8__25_), .S(SUMB_8__25_) );
  FA_X1 S2_8_26 ( .A(ab_8__26_), .B(CARRYB_7__26_), .CI(SUMB_7__27_), .CO(
        CARRYB_8__26_), .S(SUMB_8__26_) );
  FA_X1 S2_8_27 ( .A(ab_8__27_), .B(CARRYB_7__27_), .CI(SUMB_7__28_), .CO(
        CARRYB_8__27_), .S(SUMB_8__27_) );
  FA_X1 S2_8_28 ( .A(ab_8__28_), .B(CARRYB_7__28_), .CI(SUMB_7__29_), .CO(
        CARRYB_8__28_), .S(SUMB_8__28_) );
  FA_X1 S2_8_29 ( .A(ab_8__29_), .B(CARRYB_7__29_), .CI(SUMB_7__30_), .CO(
        CARRYB_8__29_), .S(SUMB_8__29_) );
  FA_X1 S3_8_30 ( .A(ab_8__30_), .B(CARRYB_7__30_), .CI(ab_7__31_), .CO(
        CARRYB_8__30_), .S(SUMB_8__30_) );
  FA_X1 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(A1_5_) );
  FA_X1 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FA_X1 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FA_X1 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FA_X1 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  FA_X1 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  FA_X1 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  FA_X1 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  FA_X1 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  FA_X1 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  FA_X1 S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  FA_X1 S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), .CO(
        CARRYB_7__17_), .S(SUMB_7__17_) );
  FA_X1 S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), .CO(
        CARRYB_7__18_), .S(SUMB_7__18_) );
  FA_X1 S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), .CO(
        CARRYB_7__19_), .S(SUMB_7__19_) );
  FA_X1 S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), .CO(
        CARRYB_7__20_), .S(SUMB_7__20_) );
  FA_X1 S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), .CO(
        CARRYB_7__21_), .S(SUMB_7__21_) );
  FA_X1 S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), .CO(
        CARRYB_7__22_), .S(SUMB_7__22_) );
  FA_X1 S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), .CO(
        CARRYB_7__23_), .S(SUMB_7__23_) );
  FA_X1 S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .CI(SUMB_6__25_), .CO(
        CARRYB_7__24_), .S(SUMB_7__24_) );
  FA_X1 S2_7_25 ( .A(ab_7__25_), .B(CARRYB_6__25_), .CI(SUMB_6__26_), .CO(
        CARRYB_7__25_), .S(SUMB_7__25_) );
  FA_X1 S2_7_26 ( .A(ab_7__26_), .B(CARRYB_6__26_), .CI(SUMB_6__27_), .CO(
        CARRYB_7__26_), .S(SUMB_7__26_) );
  FA_X1 S2_7_27 ( .A(ab_7__27_), .B(CARRYB_6__27_), .CI(SUMB_6__28_), .CO(
        CARRYB_7__27_), .S(SUMB_7__27_) );
  FA_X1 S2_7_28 ( .A(ab_7__28_), .B(CARRYB_6__28_), .CI(SUMB_6__29_), .CO(
        CARRYB_7__28_), .S(SUMB_7__28_) );
  FA_X1 S2_7_29 ( .A(ab_7__29_), .B(CARRYB_6__29_), .CI(SUMB_6__30_), .CO(
        CARRYB_7__29_), .S(SUMB_7__29_) );
  FA_X1 S3_7_30 ( .A(ab_7__30_), .B(CARRYB_6__30_), .CI(ab_6__31_), .CO(
        CARRYB_7__30_), .S(SUMB_7__30_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FA_X1 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FA_X1 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FA_X1 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  FA_X1 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  FA_X1 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  FA_X1 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  FA_X1 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  FA_X1 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  FA_X1 S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  FA_X1 S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), .CO(
        CARRYB_6__17_), .S(SUMB_6__17_) );
  FA_X1 S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), .CO(
        CARRYB_6__18_), .S(SUMB_6__18_) );
  FA_X1 S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), .CO(
        CARRYB_6__19_), .S(SUMB_6__19_) );
  FA_X1 S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), .CO(
        CARRYB_6__20_), .S(SUMB_6__20_) );
  FA_X1 S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), .CO(
        CARRYB_6__21_), .S(SUMB_6__21_) );
  FA_X1 S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), .CO(
        CARRYB_6__22_), .S(SUMB_6__22_) );
  FA_X1 S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), .CO(
        CARRYB_6__23_), .S(SUMB_6__23_) );
  FA_X1 S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), .CO(
        CARRYB_6__24_), .S(SUMB_6__24_) );
  FA_X1 S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .CI(SUMB_5__26_), .CO(
        CARRYB_6__25_), .S(SUMB_6__25_) );
  FA_X1 S2_6_26 ( .A(ab_6__26_), .B(CARRYB_5__26_), .CI(SUMB_5__27_), .CO(
        CARRYB_6__26_), .S(SUMB_6__26_) );
  FA_X1 S2_6_27 ( .A(ab_6__27_), .B(CARRYB_5__27_), .CI(SUMB_5__28_), .CO(
        CARRYB_6__27_), .S(SUMB_6__27_) );
  FA_X1 S2_6_28 ( .A(ab_6__28_), .B(CARRYB_5__28_), .CI(SUMB_5__29_), .CO(
        CARRYB_6__28_), .S(SUMB_6__28_) );
  FA_X1 S2_6_29 ( .A(ab_6__29_), .B(CARRYB_5__29_), .CI(SUMB_5__30_), .CO(
        CARRYB_6__29_), .S(SUMB_6__29_) );
  FA_X1 S3_6_30 ( .A(ab_6__30_), .B(CARRYB_5__30_), .CI(ab_5__31_), .CO(
        CARRYB_6__30_), .S(SUMB_6__30_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FA_X1 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FA_X1 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FA_X1 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  FA_X1 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  FA_X1 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  FA_X1 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  FA_X1 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  FA_X1 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  FA_X1 S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  FA_X1 S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), .CO(
        CARRYB_5__17_), .S(SUMB_5__17_) );
  FA_X1 S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), .CO(
        CARRYB_5__18_), .S(SUMB_5__18_) );
  FA_X1 S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), .CO(
        CARRYB_5__19_), .S(SUMB_5__19_) );
  FA_X1 S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), .CO(
        CARRYB_5__20_), .S(SUMB_5__20_) );
  FA_X1 S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), .CO(
        CARRYB_5__21_), .S(SUMB_5__21_) );
  FA_X1 S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), .CO(
        CARRYB_5__22_), .S(SUMB_5__22_) );
  FA_X1 S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), .CO(
        CARRYB_5__23_), .S(SUMB_5__23_) );
  FA_X1 S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), .CO(
        CARRYB_5__24_), .S(SUMB_5__24_) );
  FA_X1 S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), .CO(
        CARRYB_5__25_), .S(SUMB_5__25_) );
  FA_X1 S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .CI(SUMB_4__27_), .CO(
        CARRYB_5__26_), .S(SUMB_5__26_) );
  FA_X1 S2_5_27 ( .A(ab_5__27_), .B(CARRYB_4__27_), .CI(SUMB_4__28_), .CO(
        CARRYB_5__27_), .S(SUMB_5__27_) );
  FA_X1 S2_5_28 ( .A(ab_5__28_), .B(CARRYB_4__28_), .CI(SUMB_4__29_), .CO(
        CARRYB_5__28_), .S(SUMB_5__28_) );
  FA_X1 S2_5_29 ( .A(ab_5__29_), .B(CARRYB_4__29_), .CI(SUMB_4__30_), .CO(
        CARRYB_5__29_), .S(SUMB_5__29_) );
  FA_X1 S3_5_30 ( .A(ab_5__30_), .B(CARRYB_4__30_), .CI(ab_4__31_), .CO(
        CARRYB_5__30_), .S(SUMB_5__30_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FA_X1 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FA_X1 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FA_X1 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  FA_X1 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  FA_X1 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  FA_X1 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  FA_X1 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  FA_X1 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  FA_X1 S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  FA_X1 S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), .CO(
        CARRYB_4__17_), .S(SUMB_4__17_) );
  FA_X1 S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), .CO(
        CARRYB_4__18_), .S(SUMB_4__18_) );
  FA_X1 S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), .CO(
        CARRYB_4__19_), .S(SUMB_4__19_) );
  FA_X1 S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), .CO(
        CARRYB_4__20_), .S(SUMB_4__20_) );
  FA_X1 S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), .CO(
        CARRYB_4__21_), .S(SUMB_4__21_) );
  FA_X1 S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), .CO(
        CARRYB_4__22_), .S(SUMB_4__22_) );
  FA_X1 S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), .CO(
        CARRYB_4__23_), .S(SUMB_4__23_) );
  FA_X1 S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), .CO(
        CARRYB_4__24_), .S(SUMB_4__24_) );
  FA_X1 S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), .CO(
        CARRYB_4__25_), .S(SUMB_4__25_) );
  FA_X1 S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), .CO(
        CARRYB_4__26_), .S(SUMB_4__26_) );
  FA_X1 S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .CI(SUMB_3__28_), .CO(
        CARRYB_4__27_), .S(SUMB_4__27_) );
  FA_X1 S2_4_28 ( .A(ab_4__28_), .B(CARRYB_3__28_), .CI(SUMB_3__29_), .CO(
        CARRYB_4__28_), .S(SUMB_4__28_) );
  FA_X1 S2_4_29 ( .A(ab_4__29_), .B(CARRYB_3__29_), .CI(SUMB_3__30_), .CO(
        CARRYB_4__29_), .S(SUMB_4__29_) );
  FA_X1 S3_4_30 ( .A(ab_4__30_), .B(CARRYB_3__30_), .CI(ab_3__31_), .CO(
        CARRYB_4__30_), .S(SUMB_4__30_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FA_X1 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FA_X1 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FA_X1 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  FA_X1 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  FA_X1 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  FA_X1 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  FA_X1 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  FA_X1 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  FA_X1 S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  FA_X1 S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), .CO(
        CARRYB_3__17_), .S(SUMB_3__17_) );
  FA_X1 S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), .CO(
        CARRYB_3__18_), .S(SUMB_3__18_) );
  FA_X1 S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), .CO(
        CARRYB_3__19_), .S(SUMB_3__19_) );
  FA_X1 S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), .CO(
        CARRYB_3__20_), .S(SUMB_3__20_) );
  FA_X1 S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), .CO(
        CARRYB_3__21_), .S(SUMB_3__21_) );
  FA_X1 S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), .CO(
        CARRYB_3__22_), .S(SUMB_3__22_) );
  FA_X1 S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), .CO(
        CARRYB_3__23_), .S(SUMB_3__23_) );
  FA_X1 S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), .CO(
        CARRYB_3__24_), .S(SUMB_3__24_) );
  FA_X1 S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), .CO(
        CARRYB_3__25_), .S(SUMB_3__25_) );
  FA_X1 S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), .CO(
        CARRYB_3__26_), .S(SUMB_3__26_) );
  FA_X1 S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), .CO(
        CARRYB_3__27_), .S(SUMB_3__27_) );
  FA_X1 S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .CI(SUMB_2__29_), .CO(
        CARRYB_3__28_), .S(SUMB_3__28_) );
  FA_X1 S2_3_29 ( .A(ab_3__29_), .B(CARRYB_2__29_), .CI(SUMB_2__30_), .CO(
        CARRYB_3__29_), .S(SUMB_3__29_) );
  FA_X1 S3_3_30 ( .A(ab_3__30_), .B(CARRYB_2__30_), .CI(ab_2__31_), .CO(
        CARRYB_3__30_), .S(SUMB_3__30_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n32), .CI(n63), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n31), .CI(n62), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n30), .CI(n61), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n29), .CI(n60), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n28), .CI(n59), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n27), .CI(n58), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S2_2_6 ( .A(ab_2__6_), .B(n26), .CI(n57), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  FA_X1 S2_2_7 ( .A(ab_2__7_), .B(n25), .CI(n56), .CO(CARRYB_2__7_), .S(
        SUMB_2__7_) );
  FA_X1 S2_2_8 ( .A(ab_2__8_), .B(n24), .CI(n55), .CO(CARRYB_2__8_), .S(
        SUMB_2__8_) );
  FA_X1 S2_2_9 ( .A(ab_2__9_), .B(n23), .CI(n54), .CO(CARRYB_2__9_), .S(
        SUMB_2__9_) );
  FA_X1 S2_2_10 ( .A(ab_2__10_), .B(n22), .CI(n53), .CO(CARRYB_2__10_), .S(
        SUMB_2__10_) );
  FA_X1 S2_2_11 ( .A(ab_2__11_), .B(n21), .CI(n52), .CO(CARRYB_2__11_), .S(
        SUMB_2__11_) );
  FA_X1 S2_2_12 ( .A(ab_2__12_), .B(n20), .CI(n51), .CO(CARRYB_2__12_), .S(
        SUMB_2__12_) );
  FA_X1 S2_2_13 ( .A(ab_2__13_), .B(n19), .CI(n50), .CO(CARRYB_2__13_), .S(
        SUMB_2__13_) );
  FA_X1 S2_2_14 ( .A(ab_2__14_), .B(n18), .CI(n49), .CO(CARRYB_2__14_), .S(
        SUMB_2__14_) );
  FA_X1 S2_2_15 ( .A(ab_2__15_), .B(n17), .CI(n48), .CO(CARRYB_2__15_), .S(
        SUMB_2__15_) );
  FA_X1 S2_2_16 ( .A(ab_2__16_), .B(n16), .CI(n47), .CO(CARRYB_2__16_), .S(
        SUMB_2__16_) );
  FA_X1 S2_2_17 ( .A(ab_2__17_), .B(n15), .CI(n46), .CO(CARRYB_2__17_), .S(
        SUMB_2__17_) );
  FA_X1 S2_2_18 ( .A(ab_2__18_), .B(n14), .CI(n45), .CO(CARRYB_2__18_), .S(
        SUMB_2__18_) );
  FA_X1 S2_2_19 ( .A(ab_2__19_), .B(n13), .CI(n44), .CO(CARRYB_2__19_), .S(
        SUMB_2__19_) );
  FA_X1 S2_2_20 ( .A(ab_2__20_), .B(n12), .CI(n43), .CO(CARRYB_2__20_), .S(
        SUMB_2__20_) );
  FA_X1 S2_2_21 ( .A(ab_2__21_), .B(n11), .CI(n42), .CO(CARRYB_2__21_), .S(
        SUMB_2__21_) );
  FA_X1 S2_2_22 ( .A(ab_2__22_), .B(n10), .CI(n41), .CO(CARRYB_2__22_), .S(
        SUMB_2__22_) );
  FA_X1 S2_2_23 ( .A(ab_2__23_), .B(n9), .CI(n40), .CO(CARRYB_2__23_), .S(
        SUMB_2__23_) );
  FA_X1 S2_2_24 ( .A(ab_2__24_), .B(n8), .CI(n39), .CO(CARRYB_2__24_), .S(
        SUMB_2__24_) );
  FA_X1 S2_2_25 ( .A(ab_2__25_), .B(n7), .CI(n38), .CO(CARRYB_2__25_), .S(
        SUMB_2__25_) );
  FA_X1 S2_2_26 ( .A(ab_2__26_), .B(n6), .CI(n37), .CO(CARRYB_2__26_), .S(
        SUMB_2__26_) );
  FA_X1 S2_2_27 ( .A(ab_2__27_), .B(n5), .CI(n36), .CO(CARRYB_2__27_), .S(
        SUMB_2__27_) );
  FA_X1 S2_2_28 ( .A(ab_2__28_), .B(n4), .CI(n35), .CO(CARRYB_2__28_), .S(
        SUMB_2__28_) );
  FA_X1 S2_2_29 ( .A(ab_2__29_), .B(n3), .CI(n34), .CO(CARRYB_2__29_), .S(
        SUMB_2__29_) );
  FA_X1 S3_2_30 ( .A(ab_2__30_), .B(n33), .CI(ab_1__31_), .CO(CARRYB_2__30_), 
        .S(SUMB_2__30_) );
  simpleMultiplier_DW01_add_0 FS_1 ( .A({n317, n115, n122, n114, n121, n113, 
        n120, n112, n103, n76, n102, n75, n101, n74, n100, n80, n99, n79, n78, 
        n104, n77, n73, n70, n65, n67, n68, n71, n98, n66, n69, n72, n81, 
        A1_29_, A1_28_, A1_27_, A1_26_, A1_25_, A1_24_, A1_23_, A1_22_, A1_21_, 
        A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, A1_13_, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, A1_4_, A1_3_, A1_2_, 
        A1_1_, A1_0_}), .B({n126, n119, n125, n118, n124, n117, n123, n116, 
        n110, n93, n109, n92, n108, n91, n107, n97, n106, n96, n95, n111, n94, 
        n90, n87, n82, n84, n85, n88, n105, n83, n86, n89, A2_30_, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[63:2]) );
  AND2_X1 U2 ( .A1(ab_0__30_), .A2(ab_1__29_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__29_), .A2(ab_1__28_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__28_), .A2(ab_1__27_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__27_), .A2(ab_1__26_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__26_), .A2(ab_1__25_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__25_), .A2(ab_1__24_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__24_), .A2(ab_1__23_), .ZN(n9) );
  AND2_X1 U9 ( .A1(ab_0__23_), .A2(ab_1__22_), .ZN(n10) );
  AND2_X1 U10 ( .A1(ab_0__22_), .A2(ab_1__21_), .ZN(n11) );
  AND2_X1 U11 ( .A1(ab_0__21_), .A2(ab_1__20_), .ZN(n12) );
  AND2_X1 U12 ( .A1(ab_0__20_), .A2(ab_1__19_), .ZN(n13) );
  AND2_X1 U13 ( .A1(ab_0__19_), .A2(ab_1__18_), .ZN(n14) );
  AND2_X1 U14 ( .A1(ab_0__18_), .A2(ab_1__17_), .ZN(n15) );
  AND2_X1 U15 ( .A1(ab_0__17_), .A2(ab_1__16_), .ZN(n16) );
  AND2_X1 U16 ( .A1(ab_0__16_), .A2(ab_1__15_), .ZN(n17) );
  AND2_X1 U17 ( .A1(ab_0__15_), .A2(ab_1__14_), .ZN(n18) );
  AND2_X1 U18 ( .A1(ab_0__14_), .A2(ab_1__13_), .ZN(n19) );
  AND2_X1 U19 ( .A1(ab_0__13_), .A2(ab_1__12_), .ZN(n20) );
  AND2_X1 U20 ( .A1(ab_0__12_), .A2(ab_1__11_), .ZN(n21) );
  AND2_X1 U21 ( .A1(ab_0__11_), .A2(ab_1__10_), .ZN(n22) );
  AND2_X1 U22 ( .A1(ab_0__10_), .A2(ab_1__9_), .ZN(n23) );
  AND2_X1 U23 ( .A1(ab_0__9_), .A2(ab_1__8_), .ZN(n24) );
  AND2_X1 U24 ( .A1(ab_0__8_), .A2(ab_1__7_), .ZN(n25) );
  AND2_X1 U25 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n26) );
  AND2_X1 U26 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n27) );
  AND2_X1 U27 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n28) );
  AND2_X1 U28 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n29) );
  AND2_X1 U29 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n30) );
  AND2_X1 U30 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n31) );
  AND2_X1 U31 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n32) );
  AND2_X1 U32 ( .A1(ab_0__31_), .A2(ab_1__30_), .ZN(n33) );
  XOR2_X1 U33 ( .A(ab_1__30_), .B(ab_0__31_), .Z(n34) );
  XOR2_X1 U34 ( .A(ab_1__29_), .B(ab_0__30_), .Z(n35) );
  XOR2_X1 U35 ( .A(ab_1__28_), .B(ab_0__29_), .Z(n36) );
  XOR2_X1 U36 ( .A(ab_1__27_), .B(ab_0__28_), .Z(n37) );
  XOR2_X1 U37 ( .A(ab_1__26_), .B(ab_0__27_), .Z(n38) );
  XOR2_X1 U38 ( .A(ab_1__25_), .B(ab_0__26_), .Z(n39) );
  XOR2_X1 U39 ( .A(ab_1__24_), .B(ab_0__25_), .Z(n40) );
  XOR2_X1 U40 ( .A(ab_1__23_), .B(ab_0__24_), .Z(n41) );
  XOR2_X1 U41 ( .A(ab_1__22_), .B(ab_0__23_), .Z(n42) );
  XOR2_X1 U42 ( .A(ab_1__21_), .B(ab_0__22_), .Z(n43) );
  XOR2_X1 U43 ( .A(ab_1__20_), .B(ab_0__21_), .Z(n44) );
  XOR2_X1 U44 ( .A(ab_1__19_), .B(ab_0__20_), .Z(n45) );
  XOR2_X1 U45 ( .A(ab_1__18_), .B(ab_0__19_), .Z(n46) );
  XOR2_X1 U46 ( .A(ab_1__17_), .B(ab_0__18_), .Z(n47) );
  XOR2_X1 U47 ( .A(ab_1__16_), .B(ab_0__17_), .Z(n48) );
  XOR2_X1 U48 ( .A(ab_1__15_), .B(ab_0__16_), .Z(n49) );
  XOR2_X1 U49 ( .A(ab_1__14_), .B(ab_0__15_), .Z(n50) );
  XOR2_X1 U50 ( .A(ab_1__13_), .B(ab_0__14_), .Z(n51) );
  XOR2_X1 U51 ( .A(ab_1__12_), .B(ab_0__13_), .Z(n52) );
  XOR2_X1 U52 ( .A(ab_1__11_), .B(ab_0__12_), .Z(n53) );
  XOR2_X1 U53 ( .A(ab_1__10_), .B(ab_0__11_), .Z(n54) );
  XOR2_X1 U54 ( .A(ab_1__9_), .B(ab_0__10_), .Z(n55) );
  XOR2_X1 U55 ( .A(ab_1__8_), .B(ab_0__9_), .Z(n56) );
  XOR2_X1 U56 ( .A(ab_1__7_), .B(ab_0__8_), .Z(n57) );
  XOR2_X1 U57 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n58) );
  XOR2_X1 U58 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n59) );
  XOR2_X1 U59 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n60) );
  XOR2_X1 U60 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n61) );
  XOR2_X1 U61 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n62) );
  XOR2_X1 U62 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n63) );
  XOR2_X1 U63 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  INV_X1 U64 ( .A(CARRYB_31__31_), .ZN(n317) );
  BUF_X1 U65 ( .A(n330), .Z(n162) );
  BUF_X1 U66 ( .A(n329), .Z(n159) );
  BUF_X1 U67 ( .A(n328), .Z(n156) );
  BUF_X1 U68 ( .A(n319), .Z(n129) );
  BUF_X1 U69 ( .A(n320), .Z(n132) );
  BUF_X1 U70 ( .A(n321), .Z(n135) );
  BUF_X1 U71 ( .A(n322), .Z(n138) );
  BUF_X1 U72 ( .A(n323), .Z(n141) );
  BUF_X1 U73 ( .A(n324), .Z(n144) );
  BUF_X1 U74 ( .A(n325), .Z(n147) );
  BUF_X1 U75 ( .A(n326), .Z(n150) );
  BUF_X1 U76 ( .A(n327), .Z(n153) );
  BUF_X1 U77 ( .A(n322), .Z(n139) );
  BUF_X1 U78 ( .A(n323), .Z(n142) );
  BUF_X1 U79 ( .A(n320), .Z(n133) );
  BUF_X1 U80 ( .A(n321), .Z(n136) );
  BUF_X1 U81 ( .A(n319), .Z(n130) );
  BUF_X1 U82 ( .A(n347), .Z(n213) );
  BUF_X1 U83 ( .A(n348), .Z(n216) );
  BUF_X1 U84 ( .A(n346), .Z(n210) );
  BUF_X1 U85 ( .A(n344), .Z(n204) );
  BUF_X1 U86 ( .A(n345), .Z(n207) );
  BUF_X1 U87 ( .A(n343), .Z(n201) );
  BUF_X1 U88 ( .A(n331), .Z(n165) );
  BUF_X1 U89 ( .A(n332), .Z(n168) );
  BUF_X1 U90 ( .A(n333), .Z(n171) );
  BUF_X1 U91 ( .A(n334), .Z(n174) );
  BUF_X1 U92 ( .A(n335), .Z(n177) );
  BUF_X1 U93 ( .A(n336), .Z(n180) );
  BUF_X1 U94 ( .A(n337), .Z(n183) );
  BUF_X1 U95 ( .A(n338), .Z(n186) );
  BUF_X1 U96 ( .A(n339), .Z(n189) );
  BUF_X1 U97 ( .A(n340), .Z(n192) );
  BUF_X1 U98 ( .A(n341), .Z(n195) );
  BUF_X1 U99 ( .A(n342), .Z(n198) );
  BUF_X1 U100 ( .A(n372), .Z(n287) );
  BUF_X1 U101 ( .A(n372), .Z(n288) );
  BUF_X1 U102 ( .A(n347), .Z(n214) );
  BUF_X1 U103 ( .A(n348), .Z(n217) );
  BUF_X1 U104 ( .A(n346), .Z(n211) );
  BUF_X1 U105 ( .A(n344), .Z(n205) );
  BUF_X1 U106 ( .A(n345), .Z(n208) );
  BUF_X1 U107 ( .A(n341), .Z(n196) );
  BUF_X1 U108 ( .A(n342), .Z(n199) );
  BUF_X1 U109 ( .A(n343), .Z(n202) );
  BUF_X1 U110 ( .A(n340), .Z(n193) );
  BUF_X1 U111 ( .A(n338), .Z(n187) );
  BUF_X1 U112 ( .A(n339), .Z(n190) );
  BUF_X1 U113 ( .A(n333), .Z(n172) );
  BUF_X1 U114 ( .A(n334), .Z(n175) );
  BUF_X1 U115 ( .A(n335), .Z(n178) );
  BUF_X1 U116 ( .A(n330), .Z(n163) );
  BUF_X1 U117 ( .A(n332), .Z(n169) );
  BUF_X1 U118 ( .A(n331), .Z(n166) );
  BUF_X1 U119 ( .A(n328), .Z(n157) );
  BUF_X1 U120 ( .A(n329), .Z(n160) );
  BUF_X1 U121 ( .A(n326), .Z(n151) );
  BUF_X1 U122 ( .A(n327), .Z(n154) );
  BUF_X1 U123 ( .A(n324), .Z(n145) );
  BUF_X1 U124 ( .A(n325), .Z(n148) );
  BUF_X1 U125 ( .A(n337), .Z(n184) );
  BUF_X1 U126 ( .A(n336), .Z(n181) );
  BUF_X1 U127 ( .A(n349), .Z(n219) );
  BUF_X1 U128 ( .A(n349), .Z(n220) );
  BUF_X1 U129 ( .A(n381), .Z(n315) );
  BUF_X1 U130 ( .A(n380), .Z(n311) );
  BUF_X1 U131 ( .A(n379), .Z(n309) );
  BUF_X1 U132 ( .A(n380), .Z(n312) );
  BUF_X1 U133 ( .A(n381), .Z(n314) );
  BUF_X1 U134 ( .A(n378), .Z(n306) );
  BUF_X1 U135 ( .A(n378), .Z(n305) );
  BUF_X1 U136 ( .A(n377), .Z(n303) );
  BUF_X1 U137 ( .A(n377), .Z(n302) );
  BUF_X1 U138 ( .A(n376), .Z(n300) );
  BUF_X1 U139 ( .A(n376), .Z(n299) );
  BUF_X1 U140 ( .A(n375), .Z(n297) );
  BUF_X1 U141 ( .A(n375), .Z(n296) );
  BUF_X1 U142 ( .A(n374), .Z(n294) );
  BUF_X1 U143 ( .A(n374), .Z(n293) );
  BUF_X1 U144 ( .A(n373), .Z(n291) );
  BUF_X1 U145 ( .A(n373), .Z(n290) );
  BUF_X1 U146 ( .A(n371), .Z(n285) );
  BUF_X1 U147 ( .A(n379), .Z(n308) );
  BUF_X1 U148 ( .A(n318), .Z(n127) );
  BUF_X1 U149 ( .A(n348), .Z(n218) );
  BUF_X1 U150 ( .A(n346), .Z(n212) );
  BUF_X1 U151 ( .A(n345), .Z(n209) );
  BUF_X1 U152 ( .A(n320), .Z(n134) );
  BUF_X1 U153 ( .A(n343), .Z(n203) );
  BUF_X1 U154 ( .A(n342), .Z(n200) );
  BUF_X1 U155 ( .A(n347), .Z(n215) );
  BUF_X1 U156 ( .A(n344), .Z(n206) );
  BUF_X1 U157 ( .A(n321), .Z(n137) );
  BUF_X1 U158 ( .A(n322), .Z(n140) );
  BUF_X1 U159 ( .A(n323), .Z(n143) );
  BUF_X1 U160 ( .A(n324), .Z(n146) );
  BUF_X1 U161 ( .A(n325), .Z(n149) );
  BUF_X1 U162 ( .A(n326), .Z(n152) );
  BUF_X1 U163 ( .A(n327), .Z(n155) );
  BUF_X1 U164 ( .A(n328), .Z(n158) );
  BUF_X1 U165 ( .A(n329), .Z(n161) );
  BUF_X1 U166 ( .A(n330), .Z(n164) );
  BUF_X1 U167 ( .A(n331), .Z(n167) );
  BUF_X1 U168 ( .A(n332), .Z(n170) );
  BUF_X1 U169 ( .A(n333), .Z(n173) );
  BUF_X1 U170 ( .A(n334), .Z(n176) );
  BUF_X1 U171 ( .A(n335), .Z(n179) );
  BUF_X1 U172 ( .A(n336), .Z(n182) );
  BUF_X1 U173 ( .A(n337), .Z(n185) );
  BUF_X1 U174 ( .A(n338), .Z(n188) );
  BUF_X1 U175 ( .A(n339), .Z(n191) );
  BUF_X1 U176 ( .A(n340), .Z(n194) );
  BUF_X1 U177 ( .A(n341), .Z(n197) );
  BUF_X1 U178 ( .A(n319), .Z(n131) );
  BUF_X1 U179 ( .A(n349), .Z(n221) );
  BUF_X1 U180 ( .A(n381), .Z(n316) );
  BUF_X1 U181 ( .A(n380), .Z(n313) );
  BUF_X1 U182 ( .A(n379), .Z(n310) );
  BUF_X1 U183 ( .A(n378), .Z(n307) );
  BUF_X1 U184 ( .A(n377), .Z(n304) );
  BUF_X1 U185 ( .A(n376), .Z(n301) );
  BUF_X1 U186 ( .A(n375), .Z(n298) );
  BUF_X1 U187 ( .A(n374), .Z(n295) );
  BUF_X1 U188 ( .A(n318), .Z(n128) );
  XOR2_X1 U189 ( .A(CARRYB_31__8_), .B(SUMB_31__9_), .Z(n65) );
  XOR2_X1 U190 ( .A(CARRYB_31__3_), .B(SUMB_31__4_), .Z(n66) );
  XOR2_X1 U191 ( .A(CARRYB_31__7_), .B(SUMB_31__8_), .Z(n67) );
  XOR2_X1 U192 ( .A(CARRYB_31__6_), .B(SUMB_31__7_), .Z(n68) );
  XOR2_X1 U193 ( .A(CARRYB_31__2_), .B(SUMB_31__3_), .Z(n69) );
  XOR2_X1 U194 ( .A(CARRYB_31__9_), .B(SUMB_31__10_), .Z(n70) );
  XOR2_X1 U195 ( .A(CARRYB_31__5_), .B(SUMB_31__6_), .Z(n71) );
  XOR2_X1 U196 ( .A(CARRYB_31__1_), .B(SUMB_31__2_), .Z(n72) );
  XOR2_X1 U197 ( .A(CARRYB_31__10_), .B(SUMB_31__11_), .Z(n73) );
  XOR2_X1 U198 ( .A(CARRYB_31__18_), .B(SUMB_31__19_), .Z(n74) );
  XOR2_X1 U199 ( .A(CARRYB_31__20_), .B(SUMB_31__21_), .Z(n75) );
  XOR2_X1 U200 ( .A(CARRYB_31__22_), .B(SUMB_31__23_), .Z(n76) );
  XOR2_X1 U201 ( .A(CARRYB_31__11_), .B(SUMB_31__12_), .Z(n77) );
  XOR2_X1 U202 ( .A(CARRYB_31__13_), .B(SUMB_31__14_), .Z(n78) );
  XOR2_X1 U203 ( .A(CARRYB_31__14_), .B(SUMB_31__15_), .Z(n79) );
  XOR2_X1 U204 ( .A(CARRYB_31__16_), .B(SUMB_31__17_), .Z(n80) );
  XOR2_X1 U205 ( .A(CARRYB_31__0_), .B(SUMB_31__1_), .Z(n81) );
  AND2_X1 U206 ( .A1(CARRYB_31__7_), .A2(SUMB_31__8_), .ZN(n82) );
  AND2_X1 U207 ( .A1(CARRYB_31__2_), .A2(SUMB_31__3_), .ZN(n83) );
  AND2_X1 U208 ( .A1(CARRYB_31__6_), .A2(SUMB_31__7_), .ZN(n84) );
  AND2_X1 U209 ( .A1(CARRYB_31__5_), .A2(SUMB_31__6_), .ZN(n85) );
  AND2_X1 U210 ( .A1(CARRYB_31__1_), .A2(SUMB_31__2_), .ZN(n86) );
  AND2_X1 U211 ( .A1(CARRYB_31__8_), .A2(SUMB_31__9_), .ZN(n87) );
  AND2_X1 U212 ( .A1(CARRYB_31__4_), .A2(SUMB_31__5_), .ZN(n88) );
  AND2_X1 U213 ( .A1(CARRYB_31__0_), .A2(SUMB_31__1_), .ZN(n89) );
  AND2_X1 U214 ( .A1(CARRYB_31__9_), .A2(SUMB_31__10_), .ZN(n90) );
  AND2_X1 U215 ( .A1(CARRYB_31__17_), .A2(SUMB_31__18_), .ZN(n91) );
  AND2_X1 U216 ( .A1(CARRYB_31__19_), .A2(SUMB_31__20_), .ZN(n92) );
  AND2_X1 U217 ( .A1(CARRYB_31__21_), .A2(SUMB_31__22_), .ZN(n93) );
  AND2_X1 U218 ( .A1(CARRYB_31__10_), .A2(SUMB_31__11_), .ZN(n94) );
  AND2_X1 U219 ( .A1(CARRYB_31__12_), .A2(SUMB_31__13_), .ZN(n95) );
  AND2_X1 U220 ( .A1(CARRYB_31__13_), .A2(SUMB_31__14_), .ZN(n96) );
  AND2_X1 U221 ( .A1(CARRYB_31__15_), .A2(SUMB_31__16_), .ZN(n97) );
  XOR2_X1 U222 ( .A(CARRYB_31__4_), .B(SUMB_31__5_), .Z(n98) );
  XOR2_X1 U223 ( .A(CARRYB_31__15_), .B(SUMB_31__16_), .Z(n99) );
  XOR2_X1 U224 ( .A(CARRYB_31__17_), .B(SUMB_31__18_), .Z(n100) );
  XOR2_X1 U225 ( .A(CARRYB_31__19_), .B(SUMB_31__20_), .Z(n101) );
  XOR2_X1 U226 ( .A(CARRYB_31__21_), .B(SUMB_31__22_), .Z(n102) );
  XOR2_X1 U227 ( .A(CARRYB_31__23_), .B(SUMB_31__24_), .Z(n103) );
  XOR2_X1 U228 ( .A(CARRYB_31__12_), .B(SUMB_31__13_), .Z(n104) );
  AND2_X1 U229 ( .A1(CARRYB_31__3_), .A2(SUMB_31__4_), .ZN(n105) );
  AND2_X1 U230 ( .A1(CARRYB_31__14_), .A2(SUMB_31__15_), .ZN(n106) );
  AND2_X1 U231 ( .A1(CARRYB_31__16_), .A2(SUMB_31__17_), .ZN(n107) );
  AND2_X1 U232 ( .A1(CARRYB_31__18_), .A2(SUMB_31__19_), .ZN(n108) );
  AND2_X1 U233 ( .A1(CARRYB_31__20_), .A2(SUMB_31__21_), .ZN(n109) );
  AND2_X1 U234 ( .A1(CARRYB_31__22_), .A2(SUMB_31__23_), .ZN(n110) );
  AND2_X1 U235 ( .A1(CARRYB_31__11_), .A2(SUMB_31__12_), .ZN(n111) );
  BUF_X1 U236 ( .A(n371), .Z(n284) );
  BUF_X1 U237 ( .A(n370), .Z(n281) );
  BUF_X1 U238 ( .A(n369), .Z(n278) );
  BUF_X1 U239 ( .A(n368), .Z(n275) );
  BUF_X1 U240 ( .A(n370), .Z(n282) );
  BUF_X1 U241 ( .A(n367), .Z(n272) );
  BUF_X1 U242 ( .A(n366), .Z(n269) );
  BUF_X1 U243 ( .A(n365), .Z(n266) );
  BUF_X1 U244 ( .A(n364), .Z(n263) );
  BUF_X1 U245 ( .A(n363), .Z(n260) );
  BUF_X1 U246 ( .A(n369), .Z(n279) );
  BUF_X1 U247 ( .A(n362), .Z(n257) );
  BUF_X1 U248 ( .A(n368), .Z(n276) );
  BUF_X1 U249 ( .A(n367), .Z(n273) );
  BUF_X1 U250 ( .A(n366), .Z(n270) );
  BUF_X1 U251 ( .A(n365), .Z(n267) );
  BUF_X1 U252 ( .A(n364), .Z(n264) );
  BUF_X1 U253 ( .A(n363), .Z(n261) );
  BUF_X1 U254 ( .A(n362), .Z(n258) );
  BUF_X1 U255 ( .A(n372), .Z(n289) );
  BUF_X1 U256 ( .A(n373), .Z(n292) );
  BUF_X1 U257 ( .A(n371), .Z(n286) );
  BUF_X1 U258 ( .A(n370), .Z(n283) );
  BUF_X1 U259 ( .A(n369), .Z(n280) );
  BUF_X1 U260 ( .A(n368), .Z(n277) );
  BUF_X1 U261 ( .A(n367), .Z(n274) );
  BUF_X1 U262 ( .A(n366), .Z(n271) );
  BUF_X1 U263 ( .A(n365), .Z(n268) );
  BUF_X1 U264 ( .A(n364), .Z(n265) );
  BUF_X1 U265 ( .A(n363), .Z(n262) );
  XOR2_X1 U266 ( .A(CARRYB_31__24_), .B(SUMB_31__25_), .Z(n112) );
  XOR2_X1 U267 ( .A(CARRYB_31__26_), .B(SUMB_31__27_), .Z(n113) );
  XOR2_X1 U268 ( .A(CARRYB_31__28_), .B(SUMB_31__29_), .Z(n114) );
  XOR2_X1 U269 ( .A(CARRYB_31__30_), .B(SUMB_31__31_), .Z(n115) );
  AND2_X1 U270 ( .A1(CARRYB_31__23_), .A2(SUMB_31__24_), .ZN(n116) );
  AND2_X1 U271 ( .A1(CARRYB_31__25_), .A2(SUMB_31__26_), .ZN(n117) );
  AND2_X1 U272 ( .A1(CARRYB_31__27_), .A2(SUMB_31__28_), .ZN(n118) );
  AND2_X1 U273 ( .A1(CARRYB_31__29_), .A2(SUMB_31__30_), .ZN(n119) );
  XOR2_X1 U274 ( .A(CARRYB_31__25_), .B(SUMB_31__26_), .Z(n120) );
  XOR2_X1 U275 ( .A(CARRYB_31__27_), .B(SUMB_31__28_), .Z(n121) );
  XOR2_X1 U276 ( .A(CARRYB_31__29_), .B(SUMB_31__30_), .Z(n122) );
  AND2_X1 U277 ( .A1(CARRYB_31__24_), .A2(SUMB_31__25_), .ZN(n123) );
  AND2_X1 U278 ( .A1(CARRYB_31__26_), .A2(SUMB_31__27_), .ZN(n124) );
  AND2_X1 U279 ( .A1(CARRYB_31__28_), .A2(SUMB_31__29_), .ZN(n125) );
  AND2_X1 U280 ( .A1(CARRYB_31__30_), .A2(SUMB_31__31_), .ZN(n126) );
  BUF_X1 U281 ( .A(n361), .Z(n254) );
  BUF_X1 U282 ( .A(n360), .Z(n251) );
  BUF_X1 U283 ( .A(n359), .Z(n248) );
  BUF_X1 U284 ( .A(n358), .Z(n245) );
  BUF_X1 U285 ( .A(n357), .Z(n242) );
  BUF_X1 U286 ( .A(n356), .Z(n239) );
  BUF_X1 U287 ( .A(n355), .Z(n236) );
  BUF_X1 U288 ( .A(n354), .Z(n233) );
  BUF_X1 U289 ( .A(n353), .Z(n230) );
  BUF_X1 U290 ( .A(n361), .Z(n255) );
  BUF_X1 U291 ( .A(n360), .Z(n252) );
  BUF_X1 U292 ( .A(n359), .Z(n249) );
  BUF_X1 U293 ( .A(n358), .Z(n246) );
  BUF_X1 U294 ( .A(n357), .Z(n243) );
  BUF_X1 U295 ( .A(n356), .Z(n240) );
  BUF_X1 U296 ( .A(n355), .Z(n237) );
  BUF_X1 U297 ( .A(n354), .Z(n234) );
  BUF_X1 U298 ( .A(n362), .Z(n259) );
  BUF_X1 U299 ( .A(n361), .Z(n256) );
  BUF_X1 U300 ( .A(n360), .Z(n253) );
  BUF_X1 U301 ( .A(n359), .Z(n250) );
  BUF_X1 U302 ( .A(n358), .Z(n247) );
  BUF_X1 U303 ( .A(n357), .Z(n244) );
  BUF_X1 U304 ( .A(n356), .Z(n241) );
  BUF_X1 U305 ( .A(n355), .Z(n238) );
  BUF_X1 U306 ( .A(n354), .Z(n235) );
  BUF_X1 U307 ( .A(n353), .Z(n232) );
  BUF_X1 U308 ( .A(n352), .Z(n227) );
  BUF_X1 U309 ( .A(n351), .Z(n224) );
  BUF_X1 U310 ( .A(n350), .Z(n223) );
  BUF_X1 U311 ( .A(n353), .Z(n231) );
  BUF_X1 U312 ( .A(n352), .Z(n228) );
  BUF_X1 U313 ( .A(n351), .Z(n225) );
  BUF_X1 U314 ( .A(n350), .Z(n222) );
  BUF_X1 U315 ( .A(n352), .Z(n229) );
  BUF_X1 U316 ( .A(n351), .Z(n226) );
  INV_X1 U317 ( .A(B[31]), .ZN(n318) );
  INV_X1 U318 ( .A(A[1]), .ZN(n380) );
  INV_X1 U319 ( .A(B[30]), .ZN(n319) );
  INV_X1 U320 ( .A(B[29]), .ZN(n320) );
  INV_X1 U321 ( .A(B[28]), .ZN(n321) );
  INV_X1 U322 ( .A(B[27]), .ZN(n322) );
  INV_X1 U323 ( .A(B[26]), .ZN(n323) );
  INV_X1 U324 ( .A(B[19]), .ZN(n330) );
  INV_X1 U325 ( .A(B[20]), .ZN(n329) );
  INV_X1 U326 ( .A(A[0]), .ZN(n381) );
  INV_X1 U327 ( .A(A[2]), .ZN(n379) );
  INV_X1 U328 ( .A(B[21]), .ZN(n328) );
  INV_X1 U329 ( .A(B[25]), .ZN(n324) );
  INV_X1 U330 ( .A(B[24]), .ZN(n325) );
  INV_X1 U331 ( .A(B[23]), .ZN(n326) );
  INV_X1 U332 ( .A(B[22]), .ZN(n327) );
  INV_X1 U333 ( .A(B[2]), .ZN(n347) );
  INV_X1 U334 ( .A(B[1]), .ZN(n348) );
  INV_X1 U335 ( .A(B[3]), .ZN(n346) );
  INV_X1 U336 ( .A(B[5]), .ZN(n344) );
  INV_X1 U337 ( .A(B[4]), .ZN(n345) );
  INV_X1 U338 ( .A(B[6]), .ZN(n343) );
  INV_X1 U339 ( .A(B[18]), .ZN(n331) );
  INV_X1 U340 ( .A(B[17]), .ZN(n332) );
  INV_X1 U341 ( .A(B[16]), .ZN(n333) );
  INV_X1 U342 ( .A(B[15]), .ZN(n334) );
  INV_X1 U343 ( .A(B[14]), .ZN(n335) );
  INV_X1 U344 ( .A(B[13]), .ZN(n336) );
  INV_X1 U345 ( .A(B[12]), .ZN(n337) );
  INV_X1 U346 ( .A(B[11]), .ZN(n338) );
  INV_X1 U347 ( .A(B[10]), .ZN(n339) );
  INV_X1 U348 ( .A(B[9]), .ZN(n340) );
  INV_X1 U349 ( .A(B[8]), .ZN(n341) );
  INV_X1 U350 ( .A(B[7]), .ZN(n342) );
  INV_X1 U351 ( .A(A[3]), .ZN(n378) );
  INV_X1 U352 ( .A(A[4]), .ZN(n377) );
  INV_X1 U353 ( .A(A[5]), .ZN(n376) );
  INV_X1 U354 ( .A(A[6]), .ZN(n375) );
  INV_X1 U355 ( .A(A[7]), .ZN(n374) );
  INV_X1 U356 ( .A(A[8]), .ZN(n373) );
  INV_X1 U357 ( .A(A[9]), .ZN(n372) );
  INV_X1 U358 ( .A(A[10]), .ZN(n371) );
  INV_X1 U359 ( .A(B[0]), .ZN(n349) );
  INV_X1 U360 ( .A(A[11]), .ZN(n370) );
  INV_X1 U361 ( .A(A[12]), .ZN(n369) );
  INV_X1 U362 ( .A(A[13]), .ZN(n368) );
  INV_X1 U363 ( .A(A[14]), .ZN(n367) );
  INV_X1 U364 ( .A(A[15]), .ZN(n366) );
  INV_X1 U365 ( .A(A[16]), .ZN(n365) );
  INV_X1 U366 ( .A(A[17]), .ZN(n364) );
  INV_X1 U367 ( .A(A[18]), .ZN(n363) );
  INV_X1 U368 ( .A(A[19]), .ZN(n362) );
  INV_X1 U369 ( .A(A[20]), .ZN(n361) );
  INV_X1 U370 ( .A(A[21]), .ZN(n360) );
  INV_X1 U371 ( .A(A[22]), .ZN(n359) );
  INV_X1 U372 ( .A(A[23]), .ZN(n358) );
  INV_X1 U373 ( .A(A[24]), .ZN(n357) );
  INV_X1 U374 ( .A(A[25]), .ZN(n356) );
  INV_X1 U375 ( .A(A[26]), .ZN(n355) );
  INV_X1 U376 ( .A(A[27]), .ZN(n354) );
  INV_X1 U377 ( .A(A[28]), .ZN(n353) );
  INV_X1 U378 ( .A(A[31]), .ZN(n350) );
  INV_X1 U379 ( .A(A[29]), .ZN(n352) );
  INV_X1 U380 ( .A(A[30]), .ZN(n351) );
  NOR2_X1 U381 ( .A1(n289), .A2(n194), .ZN(ab_9__9_) );
  NOR2_X1 U382 ( .A1(n289), .A2(n197), .ZN(ab_9__8_) );
  NOR2_X1 U383 ( .A1(n289), .A2(n200), .ZN(ab_9__7_) );
  NOR2_X1 U384 ( .A1(n289), .A2(n203), .ZN(ab_9__6_) );
  NOR2_X1 U385 ( .A1(n289), .A2(n206), .ZN(ab_9__5_) );
  NOR2_X1 U386 ( .A1(n289), .A2(n209), .ZN(ab_9__4_) );
  NOR2_X1 U387 ( .A1(n289), .A2(n212), .ZN(ab_9__3_) );
  NOR2_X1 U388 ( .A1(A[9]), .A2(n127), .ZN(ab_9__31_) );
  NOR2_X1 U389 ( .A1(n288), .A2(n131), .ZN(ab_9__30_) );
  NOR2_X1 U390 ( .A1(n288), .A2(n215), .ZN(ab_9__2_) );
  NOR2_X1 U391 ( .A1(n288), .A2(n134), .ZN(ab_9__29_) );
  NOR2_X1 U392 ( .A1(n288), .A2(n137), .ZN(ab_9__28_) );
  NOR2_X1 U393 ( .A1(n288), .A2(n140), .ZN(ab_9__27_) );
  NOR2_X1 U394 ( .A1(n288), .A2(n143), .ZN(ab_9__26_) );
  NOR2_X1 U395 ( .A1(n288), .A2(n146), .ZN(ab_9__25_) );
  NOR2_X1 U396 ( .A1(n288), .A2(n149), .ZN(ab_9__24_) );
  NOR2_X1 U397 ( .A1(n288), .A2(n152), .ZN(ab_9__23_) );
  NOR2_X1 U398 ( .A1(n288), .A2(n155), .ZN(ab_9__22_) );
  NOR2_X1 U399 ( .A1(n288), .A2(n158), .ZN(ab_9__21_) );
  NOR2_X1 U400 ( .A1(n288), .A2(n161), .ZN(ab_9__20_) );
  NOR2_X1 U401 ( .A1(n287), .A2(n218), .ZN(ab_9__1_) );
  NOR2_X1 U402 ( .A1(n287), .A2(n164), .ZN(ab_9__19_) );
  NOR2_X1 U403 ( .A1(n287), .A2(n167), .ZN(ab_9__18_) );
  NOR2_X1 U404 ( .A1(n287), .A2(n170), .ZN(ab_9__17_) );
  NOR2_X1 U405 ( .A1(n287), .A2(n173), .ZN(ab_9__16_) );
  NOR2_X1 U406 ( .A1(n287), .A2(n176), .ZN(ab_9__15_) );
  NOR2_X1 U407 ( .A1(n287), .A2(n179), .ZN(ab_9__14_) );
  NOR2_X1 U408 ( .A1(n287), .A2(n182), .ZN(ab_9__13_) );
  NOR2_X1 U409 ( .A1(n287), .A2(n185), .ZN(ab_9__12_) );
  NOR2_X1 U410 ( .A1(n287), .A2(n188), .ZN(ab_9__11_) );
  NOR2_X1 U411 ( .A1(n287), .A2(n191), .ZN(ab_9__10_) );
  NOR2_X1 U412 ( .A1(n287), .A2(n221), .ZN(ab_9__0_) );
  NOR2_X1 U413 ( .A1(n194), .A2(n292), .ZN(ab_8__9_) );
  NOR2_X1 U414 ( .A1(n197), .A2(n292), .ZN(ab_8__8_) );
  NOR2_X1 U415 ( .A1(n200), .A2(n292), .ZN(ab_8__7_) );
  NOR2_X1 U416 ( .A1(n203), .A2(n292), .ZN(ab_8__6_) );
  NOR2_X1 U417 ( .A1(n206), .A2(n292), .ZN(ab_8__5_) );
  NOR2_X1 U418 ( .A1(n209), .A2(n292), .ZN(ab_8__4_) );
  NOR2_X1 U419 ( .A1(n212), .A2(n292), .ZN(ab_8__3_) );
  NOR2_X1 U420 ( .A1(A[8]), .A2(n128), .ZN(ab_8__31_) );
  NOR2_X1 U421 ( .A1(n131), .A2(n291), .ZN(ab_8__30_) );
  NOR2_X1 U422 ( .A1(n215), .A2(n291), .ZN(ab_8__2_) );
  NOR2_X1 U423 ( .A1(n134), .A2(n291), .ZN(ab_8__29_) );
  NOR2_X1 U424 ( .A1(n137), .A2(n291), .ZN(ab_8__28_) );
  NOR2_X1 U425 ( .A1(n140), .A2(n291), .ZN(ab_8__27_) );
  NOR2_X1 U426 ( .A1(n143), .A2(n291), .ZN(ab_8__26_) );
  NOR2_X1 U427 ( .A1(n146), .A2(n291), .ZN(ab_8__25_) );
  NOR2_X1 U428 ( .A1(n149), .A2(n291), .ZN(ab_8__24_) );
  NOR2_X1 U429 ( .A1(n152), .A2(n291), .ZN(ab_8__23_) );
  NOR2_X1 U430 ( .A1(n155), .A2(n291), .ZN(ab_8__22_) );
  NOR2_X1 U431 ( .A1(n158), .A2(n291), .ZN(ab_8__21_) );
  NOR2_X1 U432 ( .A1(n161), .A2(n291), .ZN(ab_8__20_) );
  NOR2_X1 U433 ( .A1(n218), .A2(n290), .ZN(ab_8__1_) );
  NOR2_X1 U434 ( .A1(n164), .A2(n290), .ZN(ab_8__19_) );
  NOR2_X1 U435 ( .A1(n167), .A2(n290), .ZN(ab_8__18_) );
  NOR2_X1 U436 ( .A1(n170), .A2(n290), .ZN(ab_8__17_) );
  NOR2_X1 U437 ( .A1(n173), .A2(n290), .ZN(ab_8__16_) );
  NOR2_X1 U438 ( .A1(n176), .A2(n290), .ZN(ab_8__15_) );
  NOR2_X1 U439 ( .A1(n179), .A2(n290), .ZN(ab_8__14_) );
  NOR2_X1 U440 ( .A1(n182), .A2(n290), .ZN(ab_8__13_) );
  NOR2_X1 U441 ( .A1(n185), .A2(n290), .ZN(ab_8__12_) );
  NOR2_X1 U442 ( .A1(n188), .A2(n290), .ZN(ab_8__11_) );
  NOR2_X1 U443 ( .A1(n191), .A2(n290), .ZN(ab_8__10_) );
  NOR2_X1 U444 ( .A1(n221), .A2(n290), .ZN(ab_8__0_) );
  NOR2_X1 U445 ( .A1(n194), .A2(n295), .ZN(ab_7__9_) );
  NOR2_X1 U446 ( .A1(n197), .A2(n295), .ZN(ab_7__8_) );
  NOR2_X1 U447 ( .A1(n200), .A2(n295), .ZN(ab_7__7_) );
  NOR2_X1 U448 ( .A1(n203), .A2(n295), .ZN(ab_7__6_) );
  NOR2_X1 U449 ( .A1(n206), .A2(n295), .ZN(ab_7__5_) );
  NOR2_X1 U450 ( .A1(n209), .A2(n295), .ZN(ab_7__4_) );
  NOR2_X1 U451 ( .A1(n212), .A2(n295), .ZN(ab_7__3_) );
  NOR2_X1 U452 ( .A1(A[7]), .A2(n128), .ZN(ab_7__31_) );
  NOR2_X1 U453 ( .A1(n131), .A2(n294), .ZN(ab_7__30_) );
  NOR2_X1 U454 ( .A1(n215), .A2(n294), .ZN(ab_7__2_) );
  NOR2_X1 U455 ( .A1(n134), .A2(n294), .ZN(ab_7__29_) );
  NOR2_X1 U456 ( .A1(n137), .A2(n294), .ZN(ab_7__28_) );
  NOR2_X1 U457 ( .A1(n140), .A2(n294), .ZN(ab_7__27_) );
  NOR2_X1 U458 ( .A1(n143), .A2(n294), .ZN(ab_7__26_) );
  NOR2_X1 U459 ( .A1(n146), .A2(n294), .ZN(ab_7__25_) );
  NOR2_X1 U460 ( .A1(n149), .A2(n294), .ZN(ab_7__24_) );
  NOR2_X1 U461 ( .A1(n152), .A2(n294), .ZN(ab_7__23_) );
  NOR2_X1 U462 ( .A1(n155), .A2(n294), .ZN(ab_7__22_) );
  NOR2_X1 U463 ( .A1(n158), .A2(n294), .ZN(ab_7__21_) );
  NOR2_X1 U464 ( .A1(n161), .A2(n294), .ZN(ab_7__20_) );
  NOR2_X1 U465 ( .A1(n218), .A2(n293), .ZN(ab_7__1_) );
  NOR2_X1 U466 ( .A1(n164), .A2(n293), .ZN(ab_7__19_) );
  NOR2_X1 U467 ( .A1(n167), .A2(n293), .ZN(ab_7__18_) );
  NOR2_X1 U468 ( .A1(n170), .A2(n293), .ZN(ab_7__17_) );
  NOR2_X1 U469 ( .A1(n173), .A2(n293), .ZN(ab_7__16_) );
  NOR2_X1 U470 ( .A1(n176), .A2(n293), .ZN(ab_7__15_) );
  NOR2_X1 U471 ( .A1(n179), .A2(n293), .ZN(ab_7__14_) );
  NOR2_X1 U472 ( .A1(n182), .A2(n293), .ZN(ab_7__13_) );
  NOR2_X1 U473 ( .A1(n185), .A2(n293), .ZN(ab_7__12_) );
  NOR2_X1 U474 ( .A1(n188), .A2(n293), .ZN(ab_7__11_) );
  NOR2_X1 U475 ( .A1(n191), .A2(n293), .ZN(ab_7__10_) );
  NOR2_X1 U476 ( .A1(n221), .A2(n293), .ZN(ab_7__0_) );
  NOR2_X1 U477 ( .A1(n194), .A2(n298), .ZN(ab_6__9_) );
  NOR2_X1 U478 ( .A1(n197), .A2(n298), .ZN(ab_6__8_) );
  NOR2_X1 U479 ( .A1(n200), .A2(n298), .ZN(ab_6__7_) );
  NOR2_X1 U480 ( .A1(n203), .A2(n298), .ZN(ab_6__6_) );
  NOR2_X1 U481 ( .A1(n206), .A2(n298), .ZN(ab_6__5_) );
  NOR2_X1 U482 ( .A1(n209), .A2(n298), .ZN(ab_6__4_) );
  NOR2_X1 U483 ( .A1(n212), .A2(n298), .ZN(ab_6__3_) );
  NOR2_X1 U484 ( .A1(A[6]), .A2(n128), .ZN(ab_6__31_) );
  NOR2_X1 U485 ( .A1(n131), .A2(n297), .ZN(ab_6__30_) );
  NOR2_X1 U486 ( .A1(n215), .A2(n297), .ZN(ab_6__2_) );
  NOR2_X1 U487 ( .A1(n134), .A2(n297), .ZN(ab_6__29_) );
  NOR2_X1 U488 ( .A1(n137), .A2(n297), .ZN(ab_6__28_) );
  NOR2_X1 U489 ( .A1(n140), .A2(n297), .ZN(ab_6__27_) );
  NOR2_X1 U490 ( .A1(n143), .A2(n297), .ZN(ab_6__26_) );
  NOR2_X1 U491 ( .A1(n146), .A2(n297), .ZN(ab_6__25_) );
  NOR2_X1 U492 ( .A1(n149), .A2(n297), .ZN(ab_6__24_) );
  NOR2_X1 U493 ( .A1(n152), .A2(n297), .ZN(ab_6__23_) );
  NOR2_X1 U494 ( .A1(n155), .A2(n297), .ZN(ab_6__22_) );
  NOR2_X1 U495 ( .A1(n158), .A2(n297), .ZN(ab_6__21_) );
  NOR2_X1 U496 ( .A1(n161), .A2(n297), .ZN(ab_6__20_) );
  NOR2_X1 U497 ( .A1(n218), .A2(n296), .ZN(ab_6__1_) );
  NOR2_X1 U498 ( .A1(n164), .A2(n296), .ZN(ab_6__19_) );
  NOR2_X1 U499 ( .A1(n167), .A2(n296), .ZN(ab_6__18_) );
  NOR2_X1 U500 ( .A1(n170), .A2(n296), .ZN(ab_6__17_) );
  NOR2_X1 U501 ( .A1(n173), .A2(n296), .ZN(ab_6__16_) );
  NOR2_X1 U502 ( .A1(n176), .A2(n296), .ZN(ab_6__15_) );
  NOR2_X1 U503 ( .A1(n179), .A2(n296), .ZN(ab_6__14_) );
  NOR2_X1 U504 ( .A1(n182), .A2(n296), .ZN(ab_6__13_) );
  NOR2_X1 U505 ( .A1(n185), .A2(n296), .ZN(ab_6__12_) );
  NOR2_X1 U506 ( .A1(n188), .A2(n296), .ZN(ab_6__11_) );
  NOR2_X1 U507 ( .A1(n191), .A2(n296), .ZN(ab_6__10_) );
  NOR2_X1 U508 ( .A1(n221), .A2(n296), .ZN(ab_6__0_) );
  NOR2_X1 U509 ( .A1(n194), .A2(n301), .ZN(ab_5__9_) );
  NOR2_X1 U510 ( .A1(n197), .A2(n301), .ZN(ab_5__8_) );
  NOR2_X1 U511 ( .A1(n200), .A2(n301), .ZN(ab_5__7_) );
  NOR2_X1 U512 ( .A1(n203), .A2(n301), .ZN(ab_5__6_) );
  NOR2_X1 U513 ( .A1(n206), .A2(n301), .ZN(ab_5__5_) );
  NOR2_X1 U514 ( .A1(n209), .A2(n301), .ZN(ab_5__4_) );
  NOR2_X1 U515 ( .A1(n212), .A2(n301), .ZN(ab_5__3_) );
  NOR2_X1 U516 ( .A1(A[5]), .A2(n128), .ZN(ab_5__31_) );
  NOR2_X1 U517 ( .A1(n131), .A2(n300), .ZN(ab_5__30_) );
  NOR2_X1 U518 ( .A1(n215), .A2(n300), .ZN(ab_5__2_) );
  NOR2_X1 U519 ( .A1(n134), .A2(n300), .ZN(ab_5__29_) );
  NOR2_X1 U520 ( .A1(n137), .A2(n300), .ZN(ab_5__28_) );
  NOR2_X1 U521 ( .A1(n140), .A2(n300), .ZN(ab_5__27_) );
  NOR2_X1 U522 ( .A1(n143), .A2(n300), .ZN(ab_5__26_) );
  NOR2_X1 U523 ( .A1(n146), .A2(n300), .ZN(ab_5__25_) );
  NOR2_X1 U524 ( .A1(n149), .A2(n300), .ZN(ab_5__24_) );
  NOR2_X1 U525 ( .A1(n152), .A2(n300), .ZN(ab_5__23_) );
  NOR2_X1 U526 ( .A1(n155), .A2(n300), .ZN(ab_5__22_) );
  NOR2_X1 U527 ( .A1(n158), .A2(n300), .ZN(ab_5__21_) );
  NOR2_X1 U528 ( .A1(n161), .A2(n300), .ZN(ab_5__20_) );
  NOR2_X1 U529 ( .A1(n218), .A2(n299), .ZN(ab_5__1_) );
  NOR2_X1 U530 ( .A1(n164), .A2(n299), .ZN(ab_5__19_) );
  NOR2_X1 U531 ( .A1(n167), .A2(n299), .ZN(ab_5__18_) );
  NOR2_X1 U532 ( .A1(n170), .A2(n299), .ZN(ab_5__17_) );
  NOR2_X1 U533 ( .A1(n173), .A2(n299), .ZN(ab_5__16_) );
  NOR2_X1 U534 ( .A1(n176), .A2(n299), .ZN(ab_5__15_) );
  NOR2_X1 U535 ( .A1(n179), .A2(n299), .ZN(ab_5__14_) );
  NOR2_X1 U536 ( .A1(n182), .A2(n299), .ZN(ab_5__13_) );
  NOR2_X1 U537 ( .A1(n185), .A2(n299), .ZN(ab_5__12_) );
  NOR2_X1 U538 ( .A1(n188), .A2(n299), .ZN(ab_5__11_) );
  NOR2_X1 U539 ( .A1(n191), .A2(n299), .ZN(ab_5__10_) );
  NOR2_X1 U540 ( .A1(n221), .A2(n299), .ZN(ab_5__0_) );
  NOR2_X1 U541 ( .A1(n194), .A2(n304), .ZN(ab_4__9_) );
  NOR2_X1 U542 ( .A1(n197), .A2(n304), .ZN(ab_4__8_) );
  NOR2_X1 U543 ( .A1(n200), .A2(n304), .ZN(ab_4__7_) );
  NOR2_X1 U544 ( .A1(n203), .A2(n304), .ZN(ab_4__6_) );
  NOR2_X1 U545 ( .A1(n206), .A2(n304), .ZN(ab_4__5_) );
  NOR2_X1 U546 ( .A1(n209), .A2(n304), .ZN(ab_4__4_) );
  NOR2_X1 U547 ( .A1(n212), .A2(n304), .ZN(ab_4__3_) );
  NOR2_X1 U548 ( .A1(A[4]), .A2(n128), .ZN(ab_4__31_) );
  NOR2_X1 U549 ( .A1(n131), .A2(n303), .ZN(ab_4__30_) );
  NOR2_X1 U550 ( .A1(n215), .A2(n303), .ZN(ab_4__2_) );
  NOR2_X1 U551 ( .A1(n134), .A2(n303), .ZN(ab_4__29_) );
  NOR2_X1 U552 ( .A1(n137), .A2(n303), .ZN(ab_4__28_) );
  NOR2_X1 U553 ( .A1(n140), .A2(n303), .ZN(ab_4__27_) );
  NOR2_X1 U554 ( .A1(n143), .A2(n303), .ZN(ab_4__26_) );
  NOR2_X1 U555 ( .A1(n146), .A2(n303), .ZN(ab_4__25_) );
  NOR2_X1 U556 ( .A1(n149), .A2(n303), .ZN(ab_4__24_) );
  NOR2_X1 U557 ( .A1(n152), .A2(n303), .ZN(ab_4__23_) );
  NOR2_X1 U558 ( .A1(n155), .A2(n303), .ZN(ab_4__22_) );
  NOR2_X1 U559 ( .A1(n158), .A2(n303), .ZN(ab_4__21_) );
  NOR2_X1 U560 ( .A1(n161), .A2(n303), .ZN(ab_4__20_) );
  NOR2_X1 U561 ( .A1(n218), .A2(n302), .ZN(ab_4__1_) );
  NOR2_X1 U562 ( .A1(n164), .A2(n302), .ZN(ab_4__19_) );
  NOR2_X1 U563 ( .A1(n167), .A2(n302), .ZN(ab_4__18_) );
  NOR2_X1 U564 ( .A1(n170), .A2(n302), .ZN(ab_4__17_) );
  NOR2_X1 U565 ( .A1(n173), .A2(n302), .ZN(ab_4__16_) );
  NOR2_X1 U566 ( .A1(n176), .A2(n302), .ZN(ab_4__15_) );
  NOR2_X1 U567 ( .A1(n179), .A2(n302), .ZN(ab_4__14_) );
  NOR2_X1 U568 ( .A1(n182), .A2(n302), .ZN(ab_4__13_) );
  NOR2_X1 U569 ( .A1(n185), .A2(n302), .ZN(ab_4__12_) );
  NOR2_X1 U570 ( .A1(n188), .A2(n302), .ZN(ab_4__11_) );
  NOR2_X1 U571 ( .A1(n191), .A2(n302), .ZN(ab_4__10_) );
  NOR2_X1 U572 ( .A1(n221), .A2(n302), .ZN(ab_4__0_) );
  NOR2_X1 U573 ( .A1(n194), .A2(n307), .ZN(ab_3__9_) );
  NOR2_X1 U574 ( .A1(n197), .A2(n307), .ZN(ab_3__8_) );
  NOR2_X1 U575 ( .A1(n200), .A2(n307), .ZN(ab_3__7_) );
  NOR2_X1 U576 ( .A1(n203), .A2(n307), .ZN(ab_3__6_) );
  NOR2_X1 U577 ( .A1(n206), .A2(n307), .ZN(ab_3__5_) );
  NOR2_X1 U578 ( .A1(n209), .A2(n307), .ZN(ab_3__4_) );
  NOR2_X1 U579 ( .A1(n212), .A2(n307), .ZN(ab_3__3_) );
  NOR2_X1 U580 ( .A1(A[3]), .A2(n128), .ZN(ab_3__31_) );
  NOR2_X1 U581 ( .A1(n131), .A2(n306), .ZN(ab_3__30_) );
  NOR2_X1 U582 ( .A1(n215), .A2(n306), .ZN(ab_3__2_) );
  NOR2_X1 U583 ( .A1(n134), .A2(n306), .ZN(ab_3__29_) );
  NOR2_X1 U584 ( .A1(n137), .A2(n306), .ZN(ab_3__28_) );
  NOR2_X1 U585 ( .A1(n140), .A2(n306), .ZN(ab_3__27_) );
  NOR2_X1 U586 ( .A1(n143), .A2(n306), .ZN(ab_3__26_) );
  NOR2_X1 U587 ( .A1(n146), .A2(n306), .ZN(ab_3__25_) );
  NOR2_X1 U588 ( .A1(n149), .A2(n306), .ZN(ab_3__24_) );
  NOR2_X1 U589 ( .A1(n152), .A2(n306), .ZN(ab_3__23_) );
  NOR2_X1 U590 ( .A1(n155), .A2(n306), .ZN(ab_3__22_) );
  NOR2_X1 U591 ( .A1(n158), .A2(n306), .ZN(ab_3__21_) );
  NOR2_X1 U592 ( .A1(n161), .A2(n306), .ZN(ab_3__20_) );
  NOR2_X1 U593 ( .A1(n218), .A2(n305), .ZN(ab_3__1_) );
  NOR2_X1 U594 ( .A1(n164), .A2(n305), .ZN(ab_3__19_) );
  NOR2_X1 U595 ( .A1(n167), .A2(n305), .ZN(ab_3__18_) );
  NOR2_X1 U596 ( .A1(n170), .A2(n305), .ZN(ab_3__17_) );
  NOR2_X1 U597 ( .A1(n173), .A2(n305), .ZN(ab_3__16_) );
  NOR2_X1 U598 ( .A1(n176), .A2(n305), .ZN(ab_3__15_) );
  NOR2_X1 U599 ( .A1(n179), .A2(n305), .ZN(ab_3__14_) );
  NOR2_X1 U600 ( .A1(n182), .A2(n305), .ZN(ab_3__13_) );
  NOR2_X1 U601 ( .A1(n185), .A2(n305), .ZN(ab_3__12_) );
  NOR2_X1 U602 ( .A1(n188), .A2(n305), .ZN(ab_3__11_) );
  NOR2_X1 U603 ( .A1(n191), .A2(n305), .ZN(ab_3__10_) );
  NOR2_X1 U604 ( .A1(n221), .A2(n305), .ZN(ab_3__0_) );
  NOR2_X1 U605 ( .A1(B[9]), .A2(n223), .ZN(ab_31__9_) );
  NOR2_X1 U606 ( .A1(B[8]), .A2(n223), .ZN(ab_31__8_) );
  NOR2_X1 U607 ( .A1(B[7]), .A2(n223), .ZN(ab_31__7_) );
  NOR2_X1 U608 ( .A1(B[6]), .A2(n223), .ZN(ab_31__6_) );
  NOR2_X1 U609 ( .A1(B[5]), .A2(n223), .ZN(ab_31__5_) );
  NOR2_X1 U610 ( .A1(B[4]), .A2(n223), .ZN(ab_31__4_) );
  NOR2_X1 U611 ( .A1(B[3]), .A2(n223), .ZN(ab_31__3_) );
  NOR2_X1 U612 ( .A1(n127), .A2(n223), .ZN(ab_31__31_) );
  NOR2_X1 U613 ( .A1(B[30]), .A2(n223), .ZN(ab_31__30_) );
  NOR2_X1 U614 ( .A1(B[2]), .A2(n223), .ZN(ab_31__2_) );
  NOR2_X1 U615 ( .A1(B[29]), .A2(n223), .ZN(ab_31__29_) );
  NOR2_X1 U616 ( .A1(B[28]), .A2(n223), .ZN(ab_31__28_) );
  NOR2_X1 U617 ( .A1(B[27]), .A2(n222), .ZN(ab_31__27_) );
  NOR2_X1 U618 ( .A1(B[26]), .A2(n222), .ZN(ab_31__26_) );
  NOR2_X1 U619 ( .A1(B[25]), .A2(n222), .ZN(ab_31__25_) );
  NOR2_X1 U620 ( .A1(B[24]), .A2(n222), .ZN(ab_31__24_) );
  NOR2_X1 U621 ( .A1(B[23]), .A2(n222), .ZN(ab_31__23_) );
  NOR2_X1 U622 ( .A1(B[22]), .A2(n222), .ZN(ab_31__22_) );
  NOR2_X1 U623 ( .A1(B[21]), .A2(n222), .ZN(ab_31__21_) );
  NOR2_X1 U624 ( .A1(B[20]), .A2(n222), .ZN(ab_31__20_) );
  NOR2_X1 U625 ( .A1(B[1]), .A2(n222), .ZN(ab_31__1_) );
  NOR2_X1 U626 ( .A1(B[19]), .A2(n222), .ZN(ab_31__19_) );
  NOR2_X1 U627 ( .A1(B[18]), .A2(n222), .ZN(ab_31__18_) );
  NOR2_X1 U628 ( .A1(B[17]), .A2(n222), .ZN(ab_31__17_) );
  NOR2_X1 U629 ( .A1(B[16]), .A2(n222), .ZN(ab_31__16_) );
  NOR2_X1 U630 ( .A1(B[15]), .A2(n222), .ZN(ab_31__15_) );
  NOR2_X1 U631 ( .A1(B[14]), .A2(n222), .ZN(ab_31__14_) );
  NOR2_X1 U632 ( .A1(B[13]), .A2(n222), .ZN(ab_31__13_) );
  NOR2_X1 U633 ( .A1(B[12]), .A2(n222), .ZN(ab_31__12_) );
  NOR2_X1 U634 ( .A1(B[11]), .A2(n222), .ZN(ab_31__11_) );
  NOR2_X1 U635 ( .A1(B[10]), .A2(n222), .ZN(ab_31__10_) );
  NOR2_X1 U636 ( .A1(B[0]), .A2(n222), .ZN(ab_31__0_) );
  NOR2_X1 U637 ( .A1(n193), .A2(n226), .ZN(ab_30__9_) );
  NOR2_X1 U638 ( .A1(n196), .A2(n226), .ZN(ab_30__8_) );
  NOR2_X1 U639 ( .A1(n199), .A2(n226), .ZN(ab_30__7_) );
  NOR2_X1 U640 ( .A1(n202), .A2(n226), .ZN(ab_30__6_) );
  NOR2_X1 U641 ( .A1(n205), .A2(n226), .ZN(ab_30__5_) );
  NOR2_X1 U642 ( .A1(n208), .A2(n226), .ZN(ab_30__4_) );
  NOR2_X1 U643 ( .A1(n211), .A2(n226), .ZN(ab_30__3_) );
  NOR2_X1 U644 ( .A1(A[30]), .A2(n128), .ZN(ab_30__31_) );
  NOR2_X1 U645 ( .A1(n130), .A2(n225), .ZN(ab_30__30_) );
  NOR2_X1 U646 ( .A1(n214), .A2(n225), .ZN(ab_30__2_) );
  NOR2_X1 U647 ( .A1(n133), .A2(n225), .ZN(ab_30__29_) );
  NOR2_X1 U648 ( .A1(n136), .A2(n225), .ZN(ab_30__28_) );
  NOR2_X1 U649 ( .A1(n139), .A2(n225), .ZN(ab_30__27_) );
  NOR2_X1 U650 ( .A1(n142), .A2(n225), .ZN(ab_30__26_) );
  NOR2_X1 U651 ( .A1(n145), .A2(n225), .ZN(ab_30__25_) );
  NOR2_X1 U652 ( .A1(n148), .A2(n225), .ZN(ab_30__24_) );
  NOR2_X1 U653 ( .A1(n151), .A2(n225), .ZN(ab_30__23_) );
  NOR2_X1 U654 ( .A1(n154), .A2(n225), .ZN(ab_30__22_) );
  NOR2_X1 U655 ( .A1(n157), .A2(n225), .ZN(ab_30__21_) );
  NOR2_X1 U656 ( .A1(n160), .A2(n225), .ZN(ab_30__20_) );
  NOR2_X1 U657 ( .A1(n217), .A2(n224), .ZN(ab_30__1_) );
  NOR2_X1 U658 ( .A1(n163), .A2(n224), .ZN(ab_30__19_) );
  NOR2_X1 U659 ( .A1(n166), .A2(n224), .ZN(ab_30__18_) );
  NOR2_X1 U660 ( .A1(n169), .A2(n224), .ZN(ab_30__17_) );
  NOR2_X1 U661 ( .A1(n172), .A2(n224), .ZN(ab_30__16_) );
  NOR2_X1 U662 ( .A1(n175), .A2(n224), .ZN(ab_30__15_) );
  NOR2_X1 U663 ( .A1(n178), .A2(n224), .ZN(ab_30__14_) );
  NOR2_X1 U664 ( .A1(n181), .A2(n224), .ZN(ab_30__13_) );
  NOR2_X1 U665 ( .A1(n184), .A2(n224), .ZN(ab_30__12_) );
  NOR2_X1 U666 ( .A1(n187), .A2(n224), .ZN(ab_30__11_) );
  NOR2_X1 U667 ( .A1(n190), .A2(n224), .ZN(ab_30__10_) );
  NOR2_X1 U668 ( .A1(n220), .A2(n224), .ZN(ab_30__0_) );
  NOR2_X1 U669 ( .A1(n193), .A2(n310), .ZN(ab_2__9_) );
  NOR2_X1 U670 ( .A1(n196), .A2(n310), .ZN(ab_2__8_) );
  NOR2_X1 U671 ( .A1(n199), .A2(n310), .ZN(ab_2__7_) );
  NOR2_X1 U672 ( .A1(n202), .A2(n310), .ZN(ab_2__6_) );
  NOR2_X1 U673 ( .A1(n205), .A2(n310), .ZN(ab_2__5_) );
  NOR2_X1 U674 ( .A1(n208), .A2(n310), .ZN(ab_2__4_) );
  NOR2_X1 U675 ( .A1(n211), .A2(n310), .ZN(ab_2__3_) );
  NOR2_X1 U676 ( .A1(A[2]), .A2(n128), .ZN(ab_2__31_) );
  NOR2_X1 U677 ( .A1(n130), .A2(n309), .ZN(ab_2__30_) );
  NOR2_X1 U678 ( .A1(n214), .A2(n309), .ZN(ab_2__2_) );
  NOR2_X1 U679 ( .A1(n133), .A2(n309), .ZN(ab_2__29_) );
  NOR2_X1 U680 ( .A1(n136), .A2(n309), .ZN(ab_2__28_) );
  NOR2_X1 U681 ( .A1(n139), .A2(n309), .ZN(ab_2__27_) );
  NOR2_X1 U682 ( .A1(n142), .A2(n309), .ZN(ab_2__26_) );
  NOR2_X1 U683 ( .A1(n145), .A2(n309), .ZN(ab_2__25_) );
  NOR2_X1 U684 ( .A1(n148), .A2(n309), .ZN(ab_2__24_) );
  NOR2_X1 U685 ( .A1(n151), .A2(n309), .ZN(ab_2__23_) );
  NOR2_X1 U686 ( .A1(n154), .A2(n309), .ZN(ab_2__22_) );
  NOR2_X1 U687 ( .A1(n157), .A2(n309), .ZN(ab_2__21_) );
  NOR2_X1 U688 ( .A1(n160), .A2(n309), .ZN(ab_2__20_) );
  NOR2_X1 U689 ( .A1(n217), .A2(n308), .ZN(ab_2__1_) );
  NOR2_X1 U690 ( .A1(n163), .A2(n308), .ZN(ab_2__19_) );
  NOR2_X1 U691 ( .A1(n166), .A2(n308), .ZN(ab_2__18_) );
  NOR2_X1 U692 ( .A1(n169), .A2(n308), .ZN(ab_2__17_) );
  NOR2_X1 U693 ( .A1(n172), .A2(n308), .ZN(ab_2__16_) );
  NOR2_X1 U694 ( .A1(n175), .A2(n308), .ZN(ab_2__15_) );
  NOR2_X1 U695 ( .A1(n178), .A2(n308), .ZN(ab_2__14_) );
  NOR2_X1 U696 ( .A1(n181), .A2(n308), .ZN(ab_2__13_) );
  NOR2_X1 U697 ( .A1(n184), .A2(n308), .ZN(ab_2__12_) );
  NOR2_X1 U698 ( .A1(n187), .A2(n308), .ZN(ab_2__11_) );
  NOR2_X1 U699 ( .A1(n190), .A2(n308), .ZN(ab_2__10_) );
  NOR2_X1 U700 ( .A1(n220), .A2(n308), .ZN(ab_2__0_) );
  NOR2_X1 U701 ( .A1(n193), .A2(n229), .ZN(ab_29__9_) );
  NOR2_X1 U702 ( .A1(n196), .A2(n229), .ZN(ab_29__8_) );
  NOR2_X1 U703 ( .A1(n199), .A2(n229), .ZN(ab_29__7_) );
  NOR2_X1 U704 ( .A1(n202), .A2(n229), .ZN(ab_29__6_) );
  NOR2_X1 U705 ( .A1(n205), .A2(n229), .ZN(ab_29__5_) );
  NOR2_X1 U706 ( .A1(n208), .A2(n229), .ZN(ab_29__4_) );
  NOR2_X1 U707 ( .A1(n211), .A2(n229), .ZN(ab_29__3_) );
  NOR2_X1 U708 ( .A1(A[29]), .A2(n128), .ZN(ab_29__31_) );
  NOR2_X1 U709 ( .A1(n130), .A2(n228), .ZN(ab_29__30_) );
  NOR2_X1 U710 ( .A1(n214), .A2(n228), .ZN(ab_29__2_) );
  NOR2_X1 U711 ( .A1(n133), .A2(n228), .ZN(ab_29__29_) );
  NOR2_X1 U712 ( .A1(n136), .A2(n228), .ZN(ab_29__28_) );
  NOR2_X1 U713 ( .A1(n139), .A2(n228), .ZN(ab_29__27_) );
  NOR2_X1 U714 ( .A1(n142), .A2(n228), .ZN(ab_29__26_) );
  NOR2_X1 U715 ( .A1(n145), .A2(n228), .ZN(ab_29__25_) );
  NOR2_X1 U716 ( .A1(n148), .A2(n228), .ZN(ab_29__24_) );
  NOR2_X1 U717 ( .A1(n151), .A2(n228), .ZN(ab_29__23_) );
  NOR2_X1 U718 ( .A1(n154), .A2(n228), .ZN(ab_29__22_) );
  NOR2_X1 U719 ( .A1(n157), .A2(n228), .ZN(ab_29__21_) );
  NOR2_X1 U720 ( .A1(n160), .A2(n228), .ZN(ab_29__20_) );
  NOR2_X1 U721 ( .A1(n217), .A2(n227), .ZN(ab_29__1_) );
  NOR2_X1 U722 ( .A1(n163), .A2(n227), .ZN(ab_29__19_) );
  NOR2_X1 U723 ( .A1(n166), .A2(n227), .ZN(ab_29__18_) );
  NOR2_X1 U724 ( .A1(n169), .A2(n227), .ZN(ab_29__17_) );
  NOR2_X1 U725 ( .A1(n172), .A2(n227), .ZN(ab_29__16_) );
  NOR2_X1 U726 ( .A1(n175), .A2(n227), .ZN(ab_29__15_) );
  NOR2_X1 U727 ( .A1(n178), .A2(n227), .ZN(ab_29__14_) );
  NOR2_X1 U728 ( .A1(n181), .A2(n227), .ZN(ab_29__13_) );
  NOR2_X1 U729 ( .A1(n184), .A2(n227), .ZN(ab_29__12_) );
  NOR2_X1 U730 ( .A1(n187), .A2(n227), .ZN(ab_29__11_) );
  NOR2_X1 U731 ( .A1(n190), .A2(n227), .ZN(ab_29__10_) );
  NOR2_X1 U732 ( .A1(n220), .A2(n227), .ZN(ab_29__0_) );
  NOR2_X1 U733 ( .A1(n193), .A2(n232), .ZN(ab_28__9_) );
  NOR2_X1 U734 ( .A1(n196), .A2(n232), .ZN(ab_28__8_) );
  NOR2_X1 U735 ( .A1(n199), .A2(n232), .ZN(ab_28__7_) );
  NOR2_X1 U736 ( .A1(n202), .A2(n232), .ZN(ab_28__6_) );
  NOR2_X1 U737 ( .A1(n205), .A2(n232), .ZN(ab_28__5_) );
  NOR2_X1 U738 ( .A1(n208), .A2(n232), .ZN(ab_28__4_) );
  NOR2_X1 U739 ( .A1(n211), .A2(n232), .ZN(ab_28__3_) );
  NOR2_X1 U740 ( .A1(A[28]), .A2(n128), .ZN(ab_28__31_) );
  NOR2_X1 U741 ( .A1(n130), .A2(n231), .ZN(ab_28__30_) );
  NOR2_X1 U742 ( .A1(n214), .A2(n231), .ZN(ab_28__2_) );
  NOR2_X1 U743 ( .A1(n133), .A2(n231), .ZN(ab_28__29_) );
  NOR2_X1 U744 ( .A1(n136), .A2(n231), .ZN(ab_28__28_) );
  NOR2_X1 U745 ( .A1(n139), .A2(n231), .ZN(ab_28__27_) );
  NOR2_X1 U746 ( .A1(n142), .A2(n231), .ZN(ab_28__26_) );
  NOR2_X1 U747 ( .A1(n145), .A2(n231), .ZN(ab_28__25_) );
  NOR2_X1 U748 ( .A1(n148), .A2(n231), .ZN(ab_28__24_) );
  NOR2_X1 U749 ( .A1(n151), .A2(n231), .ZN(ab_28__23_) );
  NOR2_X1 U750 ( .A1(n154), .A2(n231), .ZN(ab_28__22_) );
  NOR2_X1 U751 ( .A1(n157), .A2(n231), .ZN(ab_28__21_) );
  NOR2_X1 U752 ( .A1(n160), .A2(n231), .ZN(ab_28__20_) );
  NOR2_X1 U753 ( .A1(n217), .A2(n230), .ZN(ab_28__1_) );
  NOR2_X1 U754 ( .A1(n163), .A2(n230), .ZN(ab_28__19_) );
  NOR2_X1 U755 ( .A1(n166), .A2(n230), .ZN(ab_28__18_) );
  NOR2_X1 U756 ( .A1(n169), .A2(n230), .ZN(ab_28__17_) );
  NOR2_X1 U757 ( .A1(n172), .A2(n230), .ZN(ab_28__16_) );
  NOR2_X1 U758 ( .A1(n175), .A2(n230), .ZN(ab_28__15_) );
  NOR2_X1 U759 ( .A1(n178), .A2(n230), .ZN(ab_28__14_) );
  NOR2_X1 U760 ( .A1(n181), .A2(n230), .ZN(ab_28__13_) );
  NOR2_X1 U761 ( .A1(n184), .A2(n230), .ZN(ab_28__12_) );
  NOR2_X1 U762 ( .A1(n187), .A2(n230), .ZN(ab_28__11_) );
  NOR2_X1 U763 ( .A1(n190), .A2(n230), .ZN(ab_28__10_) );
  NOR2_X1 U764 ( .A1(n220), .A2(n230), .ZN(ab_28__0_) );
  NOR2_X1 U765 ( .A1(n193), .A2(n235), .ZN(ab_27__9_) );
  NOR2_X1 U766 ( .A1(n196), .A2(n235), .ZN(ab_27__8_) );
  NOR2_X1 U767 ( .A1(n199), .A2(n235), .ZN(ab_27__7_) );
  NOR2_X1 U768 ( .A1(n202), .A2(n235), .ZN(ab_27__6_) );
  NOR2_X1 U769 ( .A1(n205), .A2(n235), .ZN(ab_27__5_) );
  NOR2_X1 U770 ( .A1(n208), .A2(n235), .ZN(ab_27__4_) );
  NOR2_X1 U771 ( .A1(n211), .A2(n235), .ZN(ab_27__3_) );
  NOR2_X1 U772 ( .A1(A[27]), .A2(n128), .ZN(ab_27__31_) );
  NOR2_X1 U773 ( .A1(n130), .A2(n234), .ZN(ab_27__30_) );
  NOR2_X1 U774 ( .A1(n214), .A2(n234), .ZN(ab_27__2_) );
  NOR2_X1 U775 ( .A1(n133), .A2(n234), .ZN(ab_27__29_) );
  NOR2_X1 U776 ( .A1(n136), .A2(n234), .ZN(ab_27__28_) );
  NOR2_X1 U777 ( .A1(n139), .A2(n234), .ZN(ab_27__27_) );
  NOR2_X1 U778 ( .A1(n142), .A2(n234), .ZN(ab_27__26_) );
  NOR2_X1 U779 ( .A1(n145), .A2(n234), .ZN(ab_27__25_) );
  NOR2_X1 U780 ( .A1(n148), .A2(n234), .ZN(ab_27__24_) );
  NOR2_X1 U781 ( .A1(n151), .A2(n234), .ZN(ab_27__23_) );
  NOR2_X1 U782 ( .A1(n154), .A2(n234), .ZN(ab_27__22_) );
  NOR2_X1 U783 ( .A1(n157), .A2(n234), .ZN(ab_27__21_) );
  NOR2_X1 U784 ( .A1(n160), .A2(n234), .ZN(ab_27__20_) );
  NOR2_X1 U785 ( .A1(n217), .A2(n233), .ZN(ab_27__1_) );
  NOR2_X1 U786 ( .A1(n163), .A2(n233), .ZN(ab_27__19_) );
  NOR2_X1 U787 ( .A1(n166), .A2(n233), .ZN(ab_27__18_) );
  NOR2_X1 U788 ( .A1(n169), .A2(n233), .ZN(ab_27__17_) );
  NOR2_X1 U789 ( .A1(n172), .A2(n233), .ZN(ab_27__16_) );
  NOR2_X1 U790 ( .A1(n175), .A2(n233), .ZN(ab_27__15_) );
  NOR2_X1 U791 ( .A1(n178), .A2(n233), .ZN(ab_27__14_) );
  NOR2_X1 U792 ( .A1(n181), .A2(n233), .ZN(ab_27__13_) );
  NOR2_X1 U793 ( .A1(n184), .A2(n233), .ZN(ab_27__12_) );
  NOR2_X1 U794 ( .A1(n187), .A2(n233), .ZN(ab_27__11_) );
  NOR2_X1 U795 ( .A1(n190), .A2(n233), .ZN(ab_27__10_) );
  NOR2_X1 U796 ( .A1(n220), .A2(n233), .ZN(ab_27__0_) );
  NOR2_X1 U797 ( .A1(n193), .A2(n238), .ZN(ab_26__9_) );
  NOR2_X1 U798 ( .A1(n196), .A2(n238), .ZN(ab_26__8_) );
  NOR2_X1 U799 ( .A1(n199), .A2(n238), .ZN(ab_26__7_) );
  NOR2_X1 U800 ( .A1(n202), .A2(n238), .ZN(ab_26__6_) );
  NOR2_X1 U801 ( .A1(n205), .A2(n238), .ZN(ab_26__5_) );
  NOR2_X1 U802 ( .A1(n208), .A2(n238), .ZN(ab_26__4_) );
  NOR2_X1 U803 ( .A1(n211), .A2(n238), .ZN(ab_26__3_) );
  NOR2_X1 U804 ( .A1(A[26]), .A2(n128), .ZN(ab_26__31_) );
  NOR2_X1 U805 ( .A1(n130), .A2(n237), .ZN(ab_26__30_) );
  NOR2_X1 U806 ( .A1(n214), .A2(n237), .ZN(ab_26__2_) );
  NOR2_X1 U807 ( .A1(n133), .A2(n237), .ZN(ab_26__29_) );
  NOR2_X1 U808 ( .A1(n136), .A2(n237), .ZN(ab_26__28_) );
  NOR2_X1 U809 ( .A1(n139), .A2(n237), .ZN(ab_26__27_) );
  NOR2_X1 U810 ( .A1(n142), .A2(n237), .ZN(ab_26__26_) );
  NOR2_X1 U811 ( .A1(n145), .A2(n237), .ZN(ab_26__25_) );
  NOR2_X1 U812 ( .A1(n148), .A2(n237), .ZN(ab_26__24_) );
  NOR2_X1 U813 ( .A1(n151), .A2(n237), .ZN(ab_26__23_) );
  NOR2_X1 U814 ( .A1(n154), .A2(n237), .ZN(ab_26__22_) );
  NOR2_X1 U815 ( .A1(n157), .A2(n237), .ZN(ab_26__21_) );
  NOR2_X1 U816 ( .A1(n160), .A2(n237), .ZN(ab_26__20_) );
  NOR2_X1 U817 ( .A1(n217), .A2(n236), .ZN(ab_26__1_) );
  NOR2_X1 U818 ( .A1(n163), .A2(n236), .ZN(ab_26__19_) );
  NOR2_X1 U819 ( .A1(n166), .A2(n236), .ZN(ab_26__18_) );
  NOR2_X1 U820 ( .A1(n169), .A2(n236), .ZN(ab_26__17_) );
  NOR2_X1 U821 ( .A1(n172), .A2(n236), .ZN(ab_26__16_) );
  NOR2_X1 U822 ( .A1(n175), .A2(n236), .ZN(ab_26__15_) );
  NOR2_X1 U823 ( .A1(n178), .A2(n236), .ZN(ab_26__14_) );
  NOR2_X1 U824 ( .A1(n181), .A2(n236), .ZN(ab_26__13_) );
  NOR2_X1 U825 ( .A1(n184), .A2(n236), .ZN(ab_26__12_) );
  NOR2_X1 U826 ( .A1(n187), .A2(n236), .ZN(ab_26__11_) );
  NOR2_X1 U827 ( .A1(n190), .A2(n236), .ZN(ab_26__10_) );
  NOR2_X1 U828 ( .A1(n220), .A2(n236), .ZN(ab_26__0_) );
  NOR2_X1 U829 ( .A1(n193), .A2(n241), .ZN(ab_25__9_) );
  NOR2_X1 U830 ( .A1(n196), .A2(n241), .ZN(ab_25__8_) );
  NOR2_X1 U831 ( .A1(n199), .A2(n241), .ZN(ab_25__7_) );
  NOR2_X1 U832 ( .A1(n202), .A2(n241), .ZN(ab_25__6_) );
  NOR2_X1 U833 ( .A1(n205), .A2(n241), .ZN(ab_25__5_) );
  NOR2_X1 U834 ( .A1(n208), .A2(n241), .ZN(ab_25__4_) );
  NOR2_X1 U835 ( .A1(n211), .A2(n241), .ZN(ab_25__3_) );
  NOR2_X1 U836 ( .A1(A[25]), .A2(n128), .ZN(ab_25__31_) );
  NOR2_X1 U837 ( .A1(n130), .A2(n240), .ZN(ab_25__30_) );
  NOR2_X1 U838 ( .A1(n214), .A2(n240), .ZN(ab_25__2_) );
  NOR2_X1 U839 ( .A1(n133), .A2(n240), .ZN(ab_25__29_) );
  NOR2_X1 U840 ( .A1(n136), .A2(n240), .ZN(ab_25__28_) );
  NOR2_X1 U841 ( .A1(n139), .A2(n240), .ZN(ab_25__27_) );
  NOR2_X1 U842 ( .A1(n142), .A2(n240), .ZN(ab_25__26_) );
  NOR2_X1 U843 ( .A1(n145), .A2(n240), .ZN(ab_25__25_) );
  NOR2_X1 U844 ( .A1(n148), .A2(n240), .ZN(ab_25__24_) );
  NOR2_X1 U845 ( .A1(n151), .A2(n240), .ZN(ab_25__23_) );
  NOR2_X1 U846 ( .A1(n154), .A2(n240), .ZN(ab_25__22_) );
  NOR2_X1 U847 ( .A1(n157), .A2(n240), .ZN(ab_25__21_) );
  NOR2_X1 U848 ( .A1(n160), .A2(n240), .ZN(ab_25__20_) );
  NOR2_X1 U849 ( .A1(n217), .A2(n239), .ZN(ab_25__1_) );
  NOR2_X1 U850 ( .A1(n163), .A2(n239), .ZN(ab_25__19_) );
  NOR2_X1 U851 ( .A1(n166), .A2(n239), .ZN(ab_25__18_) );
  NOR2_X1 U852 ( .A1(n169), .A2(n239), .ZN(ab_25__17_) );
  NOR2_X1 U853 ( .A1(n172), .A2(n239), .ZN(ab_25__16_) );
  NOR2_X1 U854 ( .A1(n175), .A2(n239), .ZN(ab_25__15_) );
  NOR2_X1 U855 ( .A1(n178), .A2(n239), .ZN(ab_25__14_) );
  NOR2_X1 U856 ( .A1(n181), .A2(n239), .ZN(ab_25__13_) );
  NOR2_X1 U857 ( .A1(n184), .A2(n239), .ZN(ab_25__12_) );
  NOR2_X1 U858 ( .A1(n187), .A2(n239), .ZN(ab_25__11_) );
  NOR2_X1 U859 ( .A1(n190), .A2(n239), .ZN(ab_25__10_) );
  NOR2_X1 U860 ( .A1(n220), .A2(n239), .ZN(ab_25__0_) );
  NOR2_X1 U861 ( .A1(n193), .A2(n244), .ZN(ab_24__9_) );
  NOR2_X1 U862 ( .A1(n196), .A2(n244), .ZN(ab_24__8_) );
  NOR2_X1 U863 ( .A1(n199), .A2(n244), .ZN(ab_24__7_) );
  NOR2_X1 U864 ( .A1(n202), .A2(n244), .ZN(ab_24__6_) );
  NOR2_X1 U865 ( .A1(n205), .A2(n244), .ZN(ab_24__5_) );
  NOR2_X1 U866 ( .A1(n208), .A2(n244), .ZN(ab_24__4_) );
  NOR2_X1 U867 ( .A1(n211), .A2(n244), .ZN(ab_24__3_) );
  NOR2_X1 U868 ( .A1(A[24]), .A2(n127), .ZN(ab_24__31_) );
  NOR2_X1 U869 ( .A1(n130), .A2(n243), .ZN(ab_24__30_) );
  NOR2_X1 U870 ( .A1(n214), .A2(n243), .ZN(ab_24__2_) );
  NOR2_X1 U871 ( .A1(n133), .A2(n243), .ZN(ab_24__29_) );
  NOR2_X1 U872 ( .A1(n136), .A2(n243), .ZN(ab_24__28_) );
  NOR2_X1 U873 ( .A1(n139), .A2(n243), .ZN(ab_24__27_) );
  NOR2_X1 U874 ( .A1(n142), .A2(n243), .ZN(ab_24__26_) );
  NOR2_X1 U875 ( .A1(n145), .A2(n243), .ZN(ab_24__25_) );
  NOR2_X1 U876 ( .A1(n148), .A2(n243), .ZN(ab_24__24_) );
  NOR2_X1 U877 ( .A1(n151), .A2(n243), .ZN(ab_24__23_) );
  NOR2_X1 U878 ( .A1(n154), .A2(n243), .ZN(ab_24__22_) );
  NOR2_X1 U879 ( .A1(n157), .A2(n243), .ZN(ab_24__21_) );
  NOR2_X1 U880 ( .A1(n160), .A2(n243), .ZN(ab_24__20_) );
  NOR2_X1 U881 ( .A1(n217), .A2(n242), .ZN(ab_24__1_) );
  NOR2_X1 U882 ( .A1(n163), .A2(n242), .ZN(ab_24__19_) );
  NOR2_X1 U883 ( .A1(n166), .A2(n242), .ZN(ab_24__18_) );
  NOR2_X1 U884 ( .A1(n169), .A2(n242), .ZN(ab_24__17_) );
  NOR2_X1 U885 ( .A1(n172), .A2(n242), .ZN(ab_24__16_) );
  NOR2_X1 U886 ( .A1(n175), .A2(n242), .ZN(ab_24__15_) );
  NOR2_X1 U887 ( .A1(n178), .A2(n242), .ZN(ab_24__14_) );
  NOR2_X1 U888 ( .A1(n181), .A2(n242), .ZN(ab_24__13_) );
  NOR2_X1 U889 ( .A1(n184), .A2(n242), .ZN(ab_24__12_) );
  NOR2_X1 U890 ( .A1(n187), .A2(n242), .ZN(ab_24__11_) );
  NOR2_X1 U891 ( .A1(n190), .A2(n242), .ZN(ab_24__10_) );
  NOR2_X1 U892 ( .A1(n220), .A2(n242), .ZN(ab_24__0_) );
  NOR2_X1 U893 ( .A1(n193), .A2(n247), .ZN(ab_23__9_) );
  NOR2_X1 U894 ( .A1(n196), .A2(n247), .ZN(ab_23__8_) );
  NOR2_X1 U895 ( .A1(n199), .A2(n247), .ZN(ab_23__7_) );
  NOR2_X1 U896 ( .A1(n202), .A2(n247), .ZN(ab_23__6_) );
  NOR2_X1 U897 ( .A1(n205), .A2(n247), .ZN(ab_23__5_) );
  NOR2_X1 U898 ( .A1(n208), .A2(n247), .ZN(ab_23__4_) );
  NOR2_X1 U899 ( .A1(n211), .A2(n247), .ZN(ab_23__3_) );
  NOR2_X1 U900 ( .A1(A[23]), .A2(n127), .ZN(ab_23__31_) );
  NOR2_X1 U901 ( .A1(n130), .A2(n246), .ZN(ab_23__30_) );
  NOR2_X1 U902 ( .A1(n214), .A2(n246), .ZN(ab_23__2_) );
  NOR2_X1 U903 ( .A1(n133), .A2(n246), .ZN(ab_23__29_) );
  NOR2_X1 U904 ( .A1(n136), .A2(n246), .ZN(ab_23__28_) );
  NOR2_X1 U905 ( .A1(n139), .A2(n246), .ZN(ab_23__27_) );
  NOR2_X1 U906 ( .A1(n142), .A2(n246), .ZN(ab_23__26_) );
  NOR2_X1 U907 ( .A1(n145), .A2(n246), .ZN(ab_23__25_) );
  NOR2_X1 U908 ( .A1(n148), .A2(n246), .ZN(ab_23__24_) );
  NOR2_X1 U909 ( .A1(n151), .A2(n246), .ZN(ab_23__23_) );
  NOR2_X1 U910 ( .A1(n154), .A2(n246), .ZN(ab_23__22_) );
  NOR2_X1 U911 ( .A1(n157), .A2(n246), .ZN(ab_23__21_) );
  NOR2_X1 U912 ( .A1(n160), .A2(n246), .ZN(ab_23__20_) );
  NOR2_X1 U913 ( .A1(n217), .A2(n245), .ZN(ab_23__1_) );
  NOR2_X1 U914 ( .A1(n163), .A2(n245), .ZN(ab_23__19_) );
  NOR2_X1 U915 ( .A1(n166), .A2(n245), .ZN(ab_23__18_) );
  NOR2_X1 U916 ( .A1(n169), .A2(n245), .ZN(ab_23__17_) );
  NOR2_X1 U917 ( .A1(n172), .A2(n245), .ZN(ab_23__16_) );
  NOR2_X1 U918 ( .A1(n175), .A2(n245), .ZN(ab_23__15_) );
  NOR2_X1 U919 ( .A1(n178), .A2(n245), .ZN(ab_23__14_) );
  NOR2_X1 U920 ( .A1(n181), .A2(n245), .ZN(ab_23__13_) );
  NOR2_X1 U921 ( .A1(n184), .A2(n245), .ZN(ab_23__12_) );
  NOR2_X1 U922 ( .A1(n187), .A2(n245), .ZN(ab_23__11_) );
  NOR2_X1 U923 ( .A1(n190), .A2(n245), .ZN(ab_23__10_) );
  NOR2_X1 U924 ( .A1(n220), .A2(n245), .ZN(ab_23__0_) );
  NOR2_X1 U925 ( .A1(n193), .A2(n250), .ZN(ab_22__9_) );
  NOR2_X1 U926 ( .A1(n196), .A2(n250), .ZN(ab_22__8_) );
  NOR2_X1 U927 ( .A1(n199), .A2(n250), .ZN(ab_22__7_) );
  NOR2_X1 U928 ( .A1(n202), .A2(n250), .ZN(ab_22__6_) );
  NOR2_X1 U929 ( .A1(n205), .A2(n250), .ZN(ab_22__5_) );
  NOR2_X1 U930 ( .A1(n208), .A2(n250), .ZN(ab_22__4_) );
  NOR2_X1 U931 ( .A1(n211), .A2(n250), .ZN(ab_22__3_) );
  NOR2_X1 U932 ( .A1(A[22]), .A2(n127), .ZN(ab_22__31_) );
  NOR2_X1 U933 ( .A1(n130), .A2(n249), .ZN(ab_22__30_) );
  NOR2_X1 U934 ( .A1(n214), .A2(n249), .ZN(ab_22__2_) );
  NOR2_X1 U935 ( .A1(n133), .A2(n249), .ZN(ab_22__29_) );
  NOR2_X1 U936 ( .A1(n136), .A2(n249), .ZN(ab_22__28_) );
  NOR2_X1 U937 ( .A1(n139), .A2(n249), .ZN(ab_22__27_) );
  NOR2_X1 U938 ( .A1(n142), .A2(n249), .ZN(ab_22__26_) );
  NOR2_X1 U939 ( .A1(n145), .A2(n249), .ZN(ab_22__25_) );
  NOR2_X1 U940 ( .A1(n148), .A2(n249), .ZN(ab_22__24_) );
  NOR2_X1 U941 ( .A1(n151), .A2(n249), .ZN(ab_22__23_) );
  NOR2_X1 U942 ( .A1(n154), .A2(n249), .ZN(ab_22__22_) );
  NOR2_X1 U943 ( .A1(n157), .A2(n249), .ZN(ab_22__21_) );
  NOR2_X1 U944 ( .A1(n160), .A2(n249), .ZN(ab_22__20_) );
  NOR2_X1 U945 ( .A1(n217), .A2(n248), .ZN(ab_22__1_) );
  NOR2_X1 U946 ( .A1(n163), .A2(n248), .ZN(ab_22__19_) );
  NOR2_X1 U947 ( .A1(n166), .A2(n248), .ZN(ab_22__18_) );
  NOR2_X1 U948 ( .A1(n169), .A2(n248), .ZN(ab_22__17_) );
  NOR2_X1 U949 ( .A1(n172), .A2(n248), .ZN(ab_22__16_) );
  NOR2_X1 U950 ( .A1(n175), .A2(n248), .ZN(ab_22__15_) );
  NOR2_X1 U951 ( .A1(n178), .A2(n248), .ZN(ab_22__14_) );
  NOR2_X1 U952 ( .A1(n181), .A2(n248), .ZN(ab_22__13_) );
  NOR2_X1 U953 ( .A1(n184), .A2(n248), .ZN(ab_22__12_) );
  NOR2_X1 U954 ( .A1(n187), .A2(n248), .ZN(ab_22__11_) );
  NOR2_X1 U955 ( .A1(n190), .A2(n248), .ZN(ab_22__10_) );
  NOR2_X1 U956 ( .A1(n220), .A2(n248), .ZN(ab_22__0_) );
  NOR2_X1 U957 ( .A1(n193), .A2(n253), .ZN(ab_21__9_) );
  NOR2_X1 U958 ( .A1(n196), .A2(n253), .ZN(ab_21__8_) );
  NOR2_X1 U959 ( .A1(n199), .A2(n253), .ZN(ab_21__7_) );
  NOR2_X1 U960 ( .A1(n202), .A2(n253), .ZN(ab_21__6_) );
  NOR2_X1 U961 ( .A1(n205), .A2(n253), .ZN(ab_21__5_) );
  NOR2_X1 U962 ( .A1(n208), .A2(n253), .ZN(ab_21__4_) );
  NOR2_X1 U963 ( .A1(n211), .A2(n253), .ZN(ab_21__3_) );
  NOR2_X1 U964 ( .A1(A[21]), .A2(n127), .ZN(ab_21__31_) );
  NOR2_X1 U965 ( .A1(n130), .A2(n252), .ZN(ab_21__30_) );
  NOR2_X1 U966 ( .A1(n214), .A2(n252), .ZN(ab_21__2_) );
  NOR2_X1 U967 ( .A1(n133), .A2(n252), .ZN(ab_21__29_) );
  NOR2_X1 U968 ( .A1(n136), .A2(n252), .ZN(ab_21__28_) );
  NOR2_X1 U969 ( .A1(n139), .A2(n252), .ZN(ab_21__27_) );
  NOR2_X1 U970 ( .A1(n142), .A2(n252), .ZN(ab_21__26_) );
  NOR2_X1 U971 ( .A1(n145), .A2(n252), .ZN(ab_21__25_) );
  NOR2_X1 U972 ( .A1(n148), .A2(n252), .ZN(ab_21__24_) );
  NOR2_X1 U973 ( .A1(n151), .A2(n252), .ZN(ab_21__23_) );
  NOR2_X1 U974 ( .A1(n154), .A2(n252), .ZN(ab_21__22_) );
  NOR2_X1 U975 ( .A1(n157), .A2(n252), .ZN(ab_21__21_) );
  NOR2_X1 U976 ( .A1(n160), .A2(n252), .ZN(ab_21__20_) );
  NOR2_X1 U977 ( .A1(n217), .A2(n251), .ZN(ab_21__1_) );
  NOR2_X1 U978 ( .A1(n163), .A2(n251), .ZN(ab_21__19_) );
  NOR2_X1 U979 ( .A1(n166), .A2(n251), .ZN(ab_21__18_) );
  NOR2_X1 U980 ( .A1(n169), .A2(n251), .ZN(ab_21__17_) );
  NOR2_X1 U981 ( .A1(n172), .A2(n251), .ZN(ab_21__16_) );
  NOR2_X1 U982 ( .A1(n175), .A2(n251), .ZN(ab_21__15_) );
  NOR2_X1 U983 ( .A1(n178), .A2(n251), .ZN(ab_21__14_) );
  NOR2_X1 U984 ( .A1(n181), .A2(n251), .ZN(ab_21__13_) );
  NOR2_X1 U985 ( .A1(n184), .A2(n251), .ZN(ab_21__12_) );
  NOR2_X1 U986 ( .A1(n187), .A2(n251), .ZN(ab_21__11_) );
  NOR2_X1 U987 ( .A1(n190), .A2(n251), .ZN(ab_21__10_) );
  NOR2_X1 U988 ( .A1(n220), .A2(n251), .ZN(ab_21__0_) );
  NOR2_X1 U989 ( .A1(n193), .A2(n256), .ZN(ab_20__9_) );
  NOR2_X1 U990 ( .A1(n196), .A2(n256), .ZN(ab_20__8_) );
  NOR2_X1 U991 ( .A1(n199), .A2(n256), .ZN(ab_20__7_) );
  NOR2_X1 U992 ( .A1(n202), .A2(n256), .ZN(ab_20__6_) );
  NOR2_X1 U993 ( .A1(n205), .A2(n256), .ZN(ab_20__5_) );
  NOR2_X1 U994 ( .A1(n208), .A2(n256), .ZN(ab_20__4_) );
  NOR2_X1 U995 ( .A1(n211), .A2(n256), .ZN(ab_20__3_) );
  NOR2_X1 U996 ( .A1(A[20]), .A2(n127), .ZN(ab_20__31_) );
  NOR2_X1 U997 ( .A1(n130), .A2(n255), .ZN(ab_20__30_) );
  NOR2_X1 U998 ( .A1(n214), .A2(n255), .ZN(ab_20__2_) );
  NOR2_X1 U999 ( .A1(n133), .A2(n255), .ZN(ab_20__29_) );
  NOR2_X1 U1000 ( .A1(n136), .A2(n255), .ZN(ab_20__28_) );
  NOR2_X1 U1001 ( .A1(n139), .A2(n255), .ZN(ab_20__27_) );
  NOR2_X1 U1002 ( .A1(n142), .A2(n255), .ZN(ab_20__26_) );
  NOR2_X1 U1003 ( .A1(n145), .A2(n255), .ZN(ab_20__25_) );
  NOR2_X1 U1004 ( .A1(n148), .A2(n255), .ZN(ab_20__24_) );
  NOR2_X1 U1005 ( .A1(n151), .A2(n255), .ZN(ab_20__23_) );
  NOR2_X1 U1006 ( .A1(n154), .A2(n255), .ZN(ab_20__22_) );
  NOR2_X1 U1007 ( .A1(n157), .A2(n255), .ZN(ab_20__21_) );
  NOR2_X1 U1008 ( .A1(n160), .A2(n255), .ZN(ab_20__20_) );
  NOR2_X1 U1009 ( .A1(n217), .A2(n254), .ZN(ab_20__1_) );
  NOR2_X1 U1010 ( .A1(n163), .A2(n254), .ZN(ab_20__19_) );
  NOR2_X1 U1011 ( .A1(n166), .A2(n254), .ZN(ab_20__18_) );
  NOR2_X1 U1012 ( .A1(n169), .A2(n254), .ZN(ab_20__17_) );
  NOR2_X1 U1013 ( .A1(n172), .A2(n254), .ZN(ab_20__16_) );
  NOR2_X1 U1014 ( .A1(n175), .A2(n254), .ZN(ab_20__15_) );
  NOR2_X1 U1015 ( .A1(n178), .A2(n254), .ZN(ab_20__14_) );
  NOR2_X1 U1016 ( .A1(n181), .A2(n254), .ZN(ab_20__13_) );
  NOR2_X1 U1017 ( .A1(n184), .A2(n254), .ZN(ab_20__12_) );
  NOR2_X1 U1018 ( .A1(n187), .A2(n254), .ZN(ab_20__11_) );
  NOR2_X1 U1019 ( .A1(n190), .A2(n254), .ZN(ab_20__10_) );
  NOR2_X1 U1020 ( .A1(n220), .A2(n254), .ZN(ab_20__0_) );
  NOR2_X1 U1021 ( .A1(n192), .A2(n313), .ZN(ab_1__9_) );
  NOR2_X1 U1022 ( .A1(n195), .A2(n313), .ZN(ab_1__8_) );
  NOR2_X1 U1023 ( .A1(n198), .A2(n313), .ZN(ab_1__7_) );
  NOR2_X1 U1024 ( .A1(n201), .A2(n313), .ZN(ab_1__6_) );
  NOR2_X1 U1025 ( .A1(n204), .A2(n313), .ZN(ab_1__5_) );
  NOR2_X1 U1026 ( .A1(n207), .A2(n313), .ZN(ab_1__4_) );
  NOR2_X1 U1027 ( .A1(n210), .A2(n313), .ZN(ab_1__3_) );
  NOR2_X1 U1028 ( .A1(A[1]), .A2(n127), .ZN(ab_1__31_) );
  NOR2_X1 U1029 ( .A1(n129), .A2(n312), .ZN(ab_1__30_) );
  NOR2_X1 U1030 ( .A1(n213), .A2(n312), .ZN(ab_1__2_) );
  NOR2_X1 U1031 ( .A1(n132), .A2(n312), .ZN(ab_1__29_) );
  NOR2_X1 U1032 ( .A1(n135), .A2(n312), .ZN(ab_1__28_) );
  NOR2_X1 U1033 ( .A1(n138), .A2(n312), .ZN(ab_1__27_) );
  NOR2_X1 U1034 ( .A1(n141), .A2(n312), .ZN(ab_1__26_) );
  NOR2_X1 U1035 ( .A1(n144), .A2(n312), .ZN(ab_1__25_) );
  NOR2_X1 U1036 ( .A1(n147), .A2(n312), .ZN(ab_1__24_) );
  NOR2_X1 U1037 ( .A1(n150), .A2(n312), .ZN(ab_1__23_) );
  NOR2_X1 U1038 ( .A1(n153), .A2(n312), .ZN(ab_1__22_) );
  NOR2_X1 U1039 ( .A1(n156), .A2(n312), .ZN(ab_1__21_) );
  NOR2_X1 U1040 ( .A1(n159), .A2(n312), .ZN(ab_1__20_) );
  NOR2_X1 U1041 ( .A1(n216), .A2(n311), .ZN(ab_1__1_) );
  NOR2_X1 U1042 ( .A1(n162), .A2(n311), .ZN(ab_1__19_) );
  NOR2_X1 U1043 ( .A1(n165), .A2(n311), .ZN(ab_1__18_) );
  NOR2_X1 U1044 ( .A1(n168), .A2(n311), .ZN(ab_1__17_) );
  NOR2_X1 U1045 ( .A1(n171), .A2(n311), .ZN(ab_1__16_) );
  NOR2_X1 U1046 ( .A1(n174), .A2(n311), .ZN(ab_1__15_) );
  NOR2_X1 U1047 ( .A1(n177), .A2(n311), .ZN(ab_1__14_) );
  NOR2_X1 U1048 ( .A1(n180), .A2(n311), .ZN(ab_1__13_) );
  NOR2_X1 U1049 ( .A1(n183), .A2(n311), .ZN(ab_1__12_) );
  NOR2_X1 U1050 ( .A1(n186), .A2(n311), .ZN(ab_1__11_) );
  NOR2_X1 U1051 ( .A1(n189), .A2(n311), .ZN(ab_1__10_) );
  NOR2_X1 U1052 ( .A1(n219), .A2(n311), .ZN(ab_1__0_) );
  NOR2_X1 U1053 ( .A1(n192), .A2(n259), .ZN(ab_19__9_) );
  NOR2_X1 U1054 ( .A1(n195), .A2(n259), .ZN(ab_19__8_) );
  NOR2_X1 U1055 ( .A1(n198), .A2(n259), .ZN(ab_19__7_) );
  NOR2_X1 U1056 ( .A1(n201), .A2(n259), .ZN(ab_19__6_) );
  NOR2_X1 U1057 ( .A1(n204), .A2(n259), .ZN(ab_19__5_) );
  NOR2_X1 U1058 ( .A1(n207), .A2(n259), .ZN(ab_19__4_) );
  NOR2_X1 U1059 ( .A1(n210), .A2(n259), .ZN(ab_19__3_) );
  NOR2_X1 U1060 ( .A1(A[19]), .A2(n127), .ZN(ab_19__31_) );
  NOR2_X1 U1061 ( .A1(n129), .A2(n258), .ZN(ab_19__30_) );
  NOR2_X1 U1062 ( .A1(n213), .A2(n258), .ZN(ab_19__2_) );
  NOR2_X1 U1063 ( .A1(n132), .A2(n258), .ZN(ab_19__29_) );
  NOR2_X1 U1064 ( .A1(n135), .A2(n258), .ZN(ab_19__28_) );
  NOR2_X1 U1065 ( .A1(n138), .A2(n258), .ZN(ab_19__27_) );
  NOR2_X1 U1066 ( .A1(n141), .A2(n258), .ZN(ab_19__26_) );
  NOR2_X1 U1067 ( .A1(n144), .A2(n258), .ZN(ab_19__25_) );
  NOR2_X1 U1068 ( .A1(n147), .A2(n258), .ZN(ab_19__24_) );
  NOR2_X1 U1069 ( .A1(n150), .A2(n258), .ZN(ab_19__23_) );
  NOR2_X1 U1070 ( .A1(n153), .A2(n258), .ZN(ab_19__22_) );
  NOR2_X1 U1071 ( .A1(n156), .A2(n258), .ZN(ab_19__21_) );
  NOR2_X1 U1072 ( .A1(n159), .A2(n258), .ZN(ab_19__20_) );
  NOR2_X1 U1073 ( .A1(n216), .A2(n257), .ZN(ab_19__1_) );
  NOR2_X1 U1074 ( .A1(n162), .A2(n257), .ZN(ab_19__19_) );
  NOR2_X1 U1075 ( .A1(n165), .A2(n257), .ZN(ab_19__18_) );
  NOR2_X1 U1076 ( .A1(n168), .A2(n257), .ZN(ab_19__17_) );
  NOR2_X1 U1077 ( .A1(n171), .A2(n257), .ZN(ab_19__16_) );
  NOR2_X1 U1078 ( .A1(n174), .A2(n257), .ZN(ab_19__15_) );
  NOR2_X1 U1079 ( .A1(n177), .A2(n257), .ZN(ab_19__14_) );
  NOR2_X1 U1080 ( .A1(n180), .A2(n257), .ZN(ab_19__13_) );
  NOR2_X1 U1081 ( .A1(n183), .A2(n257), .ZN(ab_19__12_) );
  NOR2_X1 U1082 ( .A1(n186), .A2(n257), .ZN(ab_19__11_) );
  NOR2_X1 U1083 ( .A1(n189), .A2(n257), .ZN(ab_19__10_) );
  NOR2_X1 U1084 ( .A1(n219), .A2(n257), .ZN(ab_19__0_) );
  NOR2_X1 U1085 ( .A1(n192), .A2(n262), .ZN(ab_18__9_) );
  NOR2_X1 U1086 ( .A1(n195), .A2(n262), .ZN(ab_18__8_) );
  NOR2_X1 U1087 ( .A1(n198), .A2(n262), .ZN(ab_18__7_) );
  NOR2_X1 U1088 ( .A1(n201), .A2(n262), .ZN(ab_18__6_) );
  NOR2_X1 U1089 ( .A1(n204), .A2(n262), .ZN(ab_18__5_) );
  NOR2_X1 U1090 ( .A1(n207), .A2(n262), .ZN(ab_18__4_) );
  NOR2_X1 U1091 ( .A1(n210), .A2(n262), .ZN(ab_18__3_) );
  NOR2_X1 U1092 ( .A1(A[18]), .A2(n127), .ZN(ab_18__31_) );
  NOR2_X1 U1093 ( .A1(n129), .A2(n261), .ZN(ab_18__30_) );
  NOR2_X1 U1094 ( .A1(n213), .A2(n261), .ZN(ab_18__2_) );
  NOR2_X1 U1095 ( .A1(n132), .A2(n261), .ZN(ab_18__29_) );
  NOR2_X1 U1096 ( .A1(n135), .A2(n261), .ZN(ab_18__28_) );
  NOR2_X1 U1097 ( .A1(n138), .A2(n261), .ZN(ab_18__27_) );
  NOR2_X1 U1098 ( .A1(n141), .A2(n261), .ZN(ab_18__26_) );
  NOR2_X1 U1099 ( .A1(n144), .A2(n261), .ZN(ab_18__25_) );
  NOR2_X1 U1100 ( .A1(n147), .A2(n261), .ZN(ab_18__24_) );
  NOR2_X1 U1101 ( .A1(n150), .A2(n261), .ZN(ab_18__23_) );
  NOR2_X1 U1102 ( .A1(n153), .A2(n261), .ZN(ab_18__22_) );
  NOR2_X1 U1103 ( .A1(n156), .A2(n261), .ZN(ab_18__21_) );
  NOR2_X1 U1104 ( .A1(n159), .A2(n261), .ZN(ab_18__20_) );
  NOR2_X1 U1105 ( .A1(n216), .A2(n260), .ZN(ab_18__1_) );
  NOR2_X1 U1106 ( .A1(n162), .A2(n260), .ZN(ab_18__19_) );
  NOR2_X1 U1107 ( .A1(n165), .A2(n260), .ZN(ab_18__18_) );
  NOR2_X1 U1108 ( .A1(n168), .A2(n260), .ZN(ab_18__17_) );
  NOR2_X1 U1109 ( .A1(n171), .A2(n260), .ZN(ab_18__16_) );
  NOR2_X1 U1110 ( .A1(n174), .A2(n260), .ZN(ab_18__15_) );
  NOR2_X1 U1111 ( .A1(n177), .A2(n260), .ZN(ab_18__14_) );
  NOR2_X1 U1112 ( .A1(n180), .A2(n260), .ZN(ab_18__13_) );
  NOR2_X1 U1113 ( .A1(n183), .A2(n260), .ZN(ab_18__12_) );
  NOR2_X1 U1114 ( .A1(n186), .A2(n260), .ZN(ab_18__11_) );
  NOR2_X1 U1115 ( .A1(n189), .A2(n260), .ZN(ab_18__10_) );
  NOR2_X1 U1116 ( .A1(n219), .A2(n260), .ZN(ab_18__0_) );
  NOR2_X1 U1117 ( .A1(n192), .A2(n265), .ZN(ab_17__9_) );
  NOR2_X1 U1118 ( .A1(n195), .A2(n265), .ZN(ab_17__8_) );
  NOR2_X1 U1119 ( .A1(n198), .A2(n265), .ZN(ab_17__7_) );
  NOR2_X1 U1120 ( .A1(n201), .A2(n265), .ZN(ab_17__6_) );
  NOR2_X1 U1121 ( .A1(n204), .A2(n265), .ZN(ab_17__5_) );
  NOR2_X1 U1122 ( .A1(n207), .A2(n265), .ZN(ab_17__4_) );
  NOR2_X1 U1123 ( .A1(n210), .A2(n265), .ZN(ab_17__3_) );
  NOR2_X1 U1124 ( .A1(A[17]), .A2(n127), .ZN(ab_17__31_) );
  NOR2_X1 U1125 ( .A1(n129), .A2(n264), .ZN(ab_17__30_) );
  NOR2_X1 U1126 ( .A1(n213), .A2(n264), .ZN(ab_17__2_) );
  NOR2_X1 U1127 ( .A1(n132), .A2(n264), .ZN(ab_17__29_) );
  NOR2_X1 U1128 ( .A1(n135), .A2(n264), .ZN(ab_17__28_) );
  NOR2_X1 U1129 ( .A1(n138), .A2(n264), .ZN(ab_17__27_) );
  NOR2_X1 U1130 ( .A1(n141), .A2(n264), .ZN(ab_17__26_) );
  NOR2_X1 U1131 ( .A1(n144), .A2(n264), .ZN(ab_17__25_) );
  NOR2_X1 U1132 ( .A1(n147), .A2(n264), .ZN(ab_17__24_) );
  NOR2_X1 U1133 ( .A1(n150), .A2(n264), .ZN(ab_17__23_) );
  NOR2_X1 U1134 ( .A1(n153), .A2(n264), .ZN(ab_17__22_) );
  NOR2_X1 U1135 ( .A1(n156), .A2(n264), .ZN(ab_17__21_) );
  NOR2_X1 U1136 ( .A1(n159), .A2(n264), .ZN(ab_17__20_) );
  NOR2_X1 U1137 ( .A1(n216), .A2(n263), .ZN(ab_17__1_) );
  NOR2_X1 U1138 ( .A1(n162), .A2(n263), .ZN(ab_17__19_) );
  NOR2_X1 U1139 ( .A1(n165), .A2(n263), .ZN(ab_17__18_) );
  NOR2_X1 U1140 ( .A1(n168), .A2(n263), .ZN(ab_17__17_) );
  NOR2_X1 U1141 ( .A1(n171), .A2(n263), .ZN(ab_17__16_) );
  NOR2_X1 U1142 ( .A1(n174), .A2(n263), .ZN(ab_17__15_) );
  NOR2_X1 U1143 ( .A1(n177), .A2(n263), .ZN(ab_17__14_) );
  NOR2_X1 U1144 ( .A1(n180), .A2(n263), .ZN(ab_17__13_) );
  NOR2_X1 U1145 ( .A1(n183), .A2(n263), .ZN(ab_17__12_) );
  NOR2_X1 U1146 ( .A1(n186), .A2(n263), .ZN(ab_17__11_) );
  NOR2_X1 U1147 ( .A1(n189), .A2(n263), .ZN(ab_17__10_) );
  NOR2_X1 U1148 ( .A1(n219), .A2(n263), .ZN(ab_17__0_) );
  NOR2_X1 U1149 ( .A1(n192), .A2(n268), .ZN(ab_16__9_) );
  NOR2_X1 U1150 ( .A1(n195), .A2(n268), .ZN(ab_16__8_) );
  NOR2_X1 U1151 ( .A1(n198), .A2(n268), .ZN(ab_16__7_) );
  NOR2_X1 U1152 ( .A1(n201), .A2(n268), .ZN(ab_16__6_) );
  NOR2_X1 U1153 ( .A1(n204), .A2(n268), .ZN(ab_16__5_) );
  NOR2_X1 U1154 ( .A1(n207), .A2(n268), .ZN(ab_16__4_) );
  NOR2_X1 U1155 ( .A1(n210), .A2(n268), .ZN(ab_16__3_) );
  NOR2_X1 U1156 ( .A1(A[16]), .A2(n127), .ZN(ab_16__31_) );
  NOR2_X1 U1157 ( .A1(n129), .A2(n267), .ZN(ab_16__30_) );
  NOR2_X1 U1158 ( .A1(n213), .A2(n267), .ZN(ab_16__2_) );
  NOR2_X1 U1159 ( .A1(n132), .A2(n267), .ZN(ab_16__29_) );
  NOR2_X1 U1160 ( .A1(n135), .A2(n267), .ZN(ab_16__28_) );
  NOR2_X1 U1161 ( .A1(n138), .A2(n267), .ZN(ab_16__27_) );
  NOR2_X1 U1162 ( .A1(n141), .A2(n267), .ZN(ab_16__26_) );
  NOR2_X1 U1163 ( .A1(n144), .A2(n267), .ZN(ab_16__25_) );
  NOR2_X1 U1164 ( .A1(n147), .A2(n267), .ZN(ab_16__24_) );
  NOR2_X1 U1165 ( .A1(n150), .A2(n267), .ZN(ab_16__23_) );
  NOR2_X1 U1166 ( .A1(n153), .A2(n267), .ZN(ab_16__22_) );
  NOR2_X1 U1167 ( .A1(n156), .A2(n267), .ZN(ab_16__21_) );
  NOR2_X1 U1168 ( .A1(n159), .A2(n267), .ZN(ab_16__20_) );
  NOR2_X1 U1169 ( .A1(n216), .A2(n266), .ZN(ab_16__1_) );
  NOR2_X1 U1170 ( .A1(n162), .A2(n266), .ZN(ab_16__19_) );
  NOR2_X1 U1171 ( .A1(n165), .A2(n266), .ZN(ab_16__18_) );
  NOR2_X1 U1172 ( .A1(n168), .A2(n266), .ZN(ab_16__17_) );
  NOR2_X1 U1173 ( .A1(n171), .A2(n266), .ZN(ab_16__16_) );
  NOR2_X1 U1174 ( .A1(n174), .A2(n266), .ZN(ab_16__15_) );
  NOR2_X1 U1175 ( .A1(n177), .A2(n266), .ZN(ab_16__14_) );
  NOR2_X1 U1176 ( .A1(n180), .A2(n266), .ZN(ab_16__13_) );
  NOR2_X1 U1177 ( .A1(n183), .A2(n266), .ZN(ab_16__12_) );
  NOR2_X1 U1178 ( .A1(n186), .A2(n266), .ZN(ab_16__11_) );
  NOR2_X1 U1179 ( .A1(n189), .A2(n266), .ZN(ab_16__10_) );
  NOR2_X1 U1180 ( .A1(n219), .A2(n266), .ZN(ab_16__0_) );
  NOR2_X1 U1181 ( .A1(n192), .A2(n271), .ZN(ab_15__9_) );
  NOR2_X1 U1182 ( .A1(n195), .A2(n271), .ZN(ab_15__8_) );
  NOR2_X1 U1183 ( .A1(n198), .A2(n271), .ZN(ab_15__7_) );
  NOR2_X1 U1184 ( .A1(n201), .A2(n271), .ZN(ab_15__6_) );
  NOR2_X1 U1185 ( .A1(n204), .A2(n271), .ZN(ab_15__5_) );
  NOR2_X1 U1186 ( .A1(n207), .A2(n271), .ZN(ab_15__4_) );
  NOR2_X1 U1187 ( .A1(n210), .A2(n271), .ZN(ab_15__3_) );
  NOR2_X1 U1188 ( .A1(A[15]), .A2(n127), .ZN(ab_15__31_) );
  NOR2_X1 U1189 ( .A1(n129), .A2(n270), .ZN(ab_15__30_) );
  NOR2_X1 U1190 ( .A1(n213), .A2(n270), .ZN(ab_15__2_) );
  NOR2_X1 U1191 ( .A1(n132), .A2(n270), .ZN(ab_15__29_) );
  NOR2_X1 U1192 ( .A1(n135), .A2(n270), .ZN(ab_15__28_) );
  NOR2_X1 U1193 ( .A1(n138), .A2(n270), .ZN(ab_15__27_) );
  NOR2_X1 U1194 ( .A1(n141), .A2(n270), .ZN(ab_15__26_) );
  NOR2_X1 U1195 ( .A1(n144), .A2(n270), .ZN(ab_15__25_) );
  NOR2_X1 U1196 ( .A1(n147), .A2(n270), .ZN(ab_15__24_) );
  NOR2_X1 U1197 ( .A1(n150), .A2(n270), .ZN(ab_15__23_) );
  NOR2_X1 U1198 ( .A1(n153), .A2(n270), .ZN(ab_15__22_) );
  NOR2_X1 U1199 ( .A1(n156), .A2(n270), .ZN(ab_15__21_) );
  NOR2_X1 U1200 ( .A1(n159), .A2(n270), .ZN(ab_15__20_) );
  NOR2_X1 U1201 ( .A1(n216), .A2(n269), .ZN(ab_15__1_) );
  NOR2_X1 U1202 ( .A1(n162), .A2(n269), .ZN(ab_15__19_) );
  NOR2_X1 U1203 ( .A1(n165), .A2(n269), .ZN(ab_15__18_) );
  NOR2_X1 U1204 ( .A1(n168), .A2(n269), .ZN(ab_15__17_) );
  NOR2_X1 U1205 ( .A1(n171), .A2(n269), .ZN(ab_15__16_) );
  NOR2_X1 U1206 ( .A1(n174), .A2(n269), .ZN(ab_15__15_) );
  NOR2_X1 U1207 ( .A1(n177), .A2(n269), .ZN(ab_15__14_) );
  NOR2_X1 U1208 ( .A1(n180), .A2(n269), .ZN(ab_15__13_) );
  NOR2_X1 U1209 ( .A1(n183), .A2(n269), .ZN(ab_15__12_) );
  NOR2_X1 U1210 ( .A1(n186), .A2(n269), .ZN(ab_15__11_) );
  NOR2_X1 U1211 ( .A1(n189), .A2(n269), .ZN(ab_15__10_) );
  NOR2_X1 U1212 ( .A1(n219), .A2(n269), .ZN(ab_15__0_) );
  NOR2_X1 U1213 ( .A1(n192), .A2(n274), .ZN(ab_14__9_) );
  NOR2_X1 U1214 ( .A1(n195), .A2(n274), .ZN(ab_14__8_) );
  NOR2_X1 U1215 ( .A1(n198), .A2(n274), .ZN(ab_14__7_) );
  NOR2_X1 U1216 ( .A1(n201), .A2(n274), .ZN(ab_14__6_) );
  NOR2_X1 U1217 ( .A1(n204), .A2(n274), .ZN(ab_14__5_) );
  NOR2_X1 U1218 ( .A1(n207), .A2(n274), .ZN(ab_14__4_) );
  NOR2_X1 U1219 ( .A1(n210), .A2(n274), .ZN(ab_14__3_) );
  NOR2_X1 U1220 ( .A1(A[14]), .A2(n127), .ZN(ab_14__31_) );
  NOR2_X1 U1221 ( .A1(n129), .A2(n273), .ZN(ab_14__30_) );
  NOR2_X1 U1222 ( .A1(n213), .A2(n273), .ZN(ab_14__2_) );
  NOR2_X1 U1223 ( .A1(n132), .A2(n273), .ZN(ab_14__29_) );
  NOR2_X1 U1224 ( .A1(n135), .A2(n273), .ZN(ab_14__28_) );
  NOR2_X1 U1225 ( .A1(n138), .A2(n273), .ZN(ab_14__27_) );
  NOR2_X1 U1226 ( .A1(n141), .A2(n273), .ZN(ab_14__26_) );
  NOR2_X1 U1227 ( .A1(n144), .A2(n273), .ZN(ab_14__25_) );
  NOR2_X1 U1228 ( .A1(n147), .A2(n273), .ZN(ab_14__24_) );
  NOR2_X1 U1229 ( .A1(n150), .A2(n273), .ZN(ab_14__23_) );
  NOR2_X1 U1230 ( .A1(n153), .A2(n273), .ZN(ab_14__22_) );
  NOR2_X1 U1231 ( .A1(n156), .A2(n273), .ZN(ab_14__21_) );
  NOR2_X1 U1232 ( .A1(n159), .A2(n273), .ZN(ab_14__20_) );
  NOR2_X1 U1233 ( .A1(n216), .A2(n272), .ZN(ab_14__1_) );
  NOR2_X1 U1234 ( .A1(n162), .A2(n272), .ZN(ab_14__19_) );
  NOR2_X1 U1235 ( .A1(n165), .A2(n272), .ZN(ab_14__18_) );
  NOR2_X1 U1236 ( .A1(n168), .A2(n272), .ZN(ab_14__17_) );
  NOR2_X1 U1237 ( .A1(n171), .A2(n272), .ZN(ab_14__16_) );
  NOR2_X1 U1238 ( .A1(n174), .A2(n272), .ZN(ab_14__15_) );
  NOR2_X1 U1239 ( .A1(n177), .A2(n272), .ZN(ab_14__14_) );
  NOR2_X1 U1240 ( .A1(n180), .A2(n272), .ZN(ab_14__13_) );
  NOR2_X1 U1241 ( .A1(n183), .A2(n272), .ZN(ab_14__12_) );
  NOR2_X1 U1242 ( .A1(n186), .A2(n272), .ZN(ab_14__11_) );
  NOR2_X1 U1243 ( .A1(n189), .A2(n272), .ZN(ab_14__10_) );
  NOR2_X1 U1244 ( .A1(n219), .A2(n272), .ZN(ab_14__0_) );
  NOR2_X1 U1245 ( .A1(n192), .A2(n277), .ZN(ab_13__9_) );
  NOR2_X1 U1246 ( .A1(n195), .A2(n277), .ZN(ab_13__8_) );
  NOR2_X1 U1247 ( .A1(n198), .A2(n277), .ZN(ab_13__7_) );
  NOR2_X1 U1248 ( .A1(n201), .A2(n277), .ZN(ab_13__6_) );
  NOR2_X1 U1249 ( .A1(n204), .A2(n277), .ZN(ab_13__5_) );
  NOR2_X1 U1250 ( .A1(n207), .A2(n277), .ZN(ab_13__4_) );
  NOR2_X1 U1251 ( .A1(n210), .A2(n277), .ZN(ab_13__3_) );
  NOR2_X1 U1252 ( .A1(A[13]), .A2(n127), .ZN(ab_13__31_) );
  NOR2_X1 U1253 ( .A1(n129), .A2(n276), .ZN(ab_13__30_) );
  NOR2_X1 U1254 ( .A1(n213), .A2(n276), .ZN(ab_13__2_) );
  NOR2_X1 U1255 ( .A1(n132), .A2(n276), .ZN(ab_13__29_) );
  NOR2_X1 U1256 ( .A1(n135), .A2(n276), .ZN(ab_13__28_) );
  NOR2_X1 U1257 ( .A1(n138), .A2(n276), .ZN(ab_13__27_) );
  NOR2_X1 U1258 ( .A1(n141), .A2(n276), .ZN(ab_13__26_) );
  NOR2_X1 U1259 ( .A1(n144), .A2(n276), .ZN(ab_13__25_) );
  NOR2_X1 U1260 ( .A1(n147), .A2(n276), .ZN(ab_13__24_) );
  NOR2_X1 U1261 ( .A1(n150), .A2(n276), .ZN(ab_13__23_) );
  NOR2_X1 U1262 ( .A1(n153), .A2(n276), .ZN(ab_13__22_) );
  NOR2_X1 U1263 ( .A1(n156), .A2(n276), .ZN(ab_13__21_) );
  NOR2_X1 U1264 ( .A1(n159), .A2(n276), .ZN(ab_13__20_) );
  NOR2_X1 U1265 ( .A1(n216), .A2(n275), .ZN(ab_13__1_) );
  NOR2_X1 U1266 ( .A1(n162), .A2(n275), .ZN(ab_13__19_) );
  NOR2_X1 U1267 ( .A1(n165), .A2(n275), .ZN(ab_13__18_) );
  NOR2_X1 U1268 ( .A1(n168), .A2(n275), .ZN(ab_13__17_) );
  NOR2_X1 U1269 ( .A1(n171), .A2(n275), .ZN(ab_13__16_) );
  NOR2_X1 U1270 ( .A1(n174), .A2(n275), .ZN(ab_13__15_) );
  NOR2_X1 U1271 ( .A1(n177), .A2(n275), .ZN(ab_13__14_) );
  NOR2_X1 U1272 ( .A1(n180), .A2(n275), .ZN(ab_13__13_) );
  NOR2_X1 U1273 ( .A1(n183), .A2(n275), .ZN(ab_13__12_) );
  NOR2_X1 U1274 ( .A1(n186), .A2(n275), .ZN(ab_13__11_) );
  NOR2_X1 U1275 ( .A1(n189), .A2(n275), .ZN(ab_13__10_) );
  NOR2_X1 U1276 ( .A1(n219), .A2(n275), .ZN(ab_13__0_) );
  NOR2_X1 U1277 ( .A1(n192), .A2(n280), .ZN(ab_12__9_) );
  NOR2_X1 U1278 ( .A1(n195), .A2(n280), .ZN(ab_12__8_) );
  NOR2_X1 U1279 ( .A1(n198), .A2(n280), .ZN(ab_12__7_) );
  NOR2_X1 U1280 ( .A1(n201), .A2(n280), .ZN(ab_12__6_) );
  NOR2_X1 U1281 ( .A1(n204), .A2(n280), .ZN(ab_12__5_) );
  NOR2_X1 U1282 ( .A1(n207), .A2(n280), .ZN(ab_12__4_) );
  NOR2_X1 U1283 ( .A1(n210), .A2(n280), .ZN(ab_12__3_) );
  NOR2_X1 U1284 ( .A1(A[12]), .A2(n127), .ZN(ab_12__31_) );
  NOR2_X1 U1285 ( .A1(n129), .A2(n279), .ZN(ab_12__30_) );
  NOR2_X1 U1286 ( .A1(n213), .A2(n279), .ZN(ab_12__2_) );
  NOR2_X1 U1287 ( .A1(n132), .A2(n279), .ZN(ab_12__29_) );
  NOR2_X1 U1288 ( .A1(n135), .A2(n279), .ZN(ab_12__28_) );
  NOR2_X1 U1289 ( .A1(n138), .A2(n279), .ZN(ab_12__27_) );
  NOR2_X1 U1290 ( .A1(n141), .A2(n279), .ZN(ab_12__26_) );
  NOR2_X1 U1291 ( .A1(n144), .A2(n279), .ZN(ab_12__25_) );
  NOR2_X1 U1292 ( .A1(n147), .A2(n279), .ZN(ab_12__24_) );
  NOR2_X1 U1293 ( .A1(n150), .A2(n279), .ZN(ab_12__23_) );
  NOR2_X1 U1294 ( .A1(n153), .A2(n279), .ZN(ab_12__22_) );
  NOR2_X1 U1295 ( .A1(n156), .A2(n279), .ZN(ab_12__21_) );
  NOR2_X1 U1296 ( .A1(n159), .A2(n279), .ZN(ab_12__20_) );
  NOR2_X1 U1297 ( .A1(n216), .A2(n278), .ZN(ab_12__1_) );
  NOR2_X1 U1298 ( .A1(n162), .A2(n278), .ZN(ab_12__19_) );
  NOR2_X1 U1299 ( .A1(n165), .A2(n278), .ZN(ab_12__18_) );
  NOR2_X1 U1300 ( .A1(n168), .A2(n278), .ZN(ab_12__17_) );
  NOR2_X1 U1301 ( .A1(n171), .A2(n278), .ZN(ab_12__16_) );
  NOR2_X1 U1302 ( .A1(n174), .A2(n278), .ZN(ab_12__15_) );
  NOR2_X1 U1303 ( .A1(n177), .A2(n278), .ZN(ab_12__14_) );
  NOR2_X1 U1304 ( .A1(n180), .A2(n278), .ZN(ab_12__13_) );
  NOR2_X1 U1305 ( .A1(n183), .A2(n278), .ZN(ab_12__12_) );
  NOR2_X1 U1306 ( .A1(n186), .A2(n278), .ZN(ab_12__11_) );
  NOR2_X1 U1307 ( .A1(n189), .A2(n278), .ZN(ab_12__10_) );
  NOR2_X1 U1308 ( .A1(n219), .A2(n278), .ZN(ab_12__0_) );
  NOR2_X1 U1309 ( .A1(n192), .A2(n283), .ZN(ab_11__9_) );
  NOR2_X1 U1310 ( .A1(n195), .A2(n283), .ZN(ab_11__8_) );
  NOR2_X1 U1311 ( .A1(n198), .A2(n283), .ZN(ab_11__7_) );
  NOR2_X1 U1312 ( .A1(n201), .A2(n283), .ZN(ab_11__6_) );
  NOR2_X1 U1313 ( .A1(n204), .A2(n283), .ZN(ab_11__5_) );
  NOR2_X1 U1314 ( .A1(n207), .A2(n283), .ZN(ab_11__4_) );
  NOR2_X1 U1315 ( .A1(n210), .A2(n283), .ZN(ab_11__3_) );
  NOR2_X1 U1316 ( .A1(A[11]), .A2(n127), .ZN(ab_11__31_) );
  NOR2_X1 U1317 ( .A1(n129), .A2(n282), .ZN(ab_11__30_) );
  NOR2_X1 U1318 ( .A1(n213), .A2(n282), .ZN(ab_11__2_) );
  NOR2_X1 U1319 ( .A1(n132), .A2(n282), .ZN(ab_11__29_) );
  NOR2_X1 U1320 ( .A1(n135), .A2(n282), .ZN(ab_11__28_) );
  NOR2_X1 U1321 ( .A1(n138), .A2(n282), .ZN(ab_11__27_) );
  NOR2_X1 U1322 ( .A1(n141), .A2(n282), .ZN(ab_11__26_) );
  NOR2_X1 U1323 ( .A1(n144), .A2(n282), .ZN(ab_11__25_) );
  NOR2_X1 U1324 ( .A1(n147), .A2(n282), .ZN(ab_11__24_) );
  NOR2_X1 U1325 ( .A1(n150), .A2(n282), .ZN(ab_11__23_) );
  NOR2_X1 U1326 ( .A1(n153), .A2(n282), .ZN(ab_11__22_) );
  NOR2_X1 U1327 ( .A1(n156), .A2(n282), .ZN(ab_11__21_) );
  NOR2_X1 U1328 ( .A1(n159), .A2(n282), .ZN(ab_11__20_) );
  NOR2_X1 U1329 ( .A1(n216), .A2(n281), .ZN(ab_11__1_) );
  NOR2_X1 U1330 ( .A1(n162), .A2(n281), .ZN(ab_11__19_) );
  NOR2_X1 U1331 ( .A1(n165), .A2(n281), .ZN(ab_11__18_) );
  NOR2_X1 U1332 ( .A1(n168), .A2(n281), .ZN(ab_11__17_) );
  NOR2_X1 U1333 ( .A1(n171), .A2(n281), .ZN(ab_11__16_) );
  NOR2_X1 U1334 ( .A1(n174), .A2(n281), .ZN(ab_11__15_) );
  NOR2_X1 U1335 ( .A1(n177), .A2(n281), .ZN(ab_11__14_) );
  NOR2_X1 U1336 ( .A1(n180), .A2(n281), .ZN(ab_11__13_) );
  NOR2_X1 U1337 ( .A1(n183), .A2(n281), .ZN(ab_11__12_) );
  NOR2_X1 U1338 ( .A1(n186), .A2(n281), .ZN(ab_11__11_) );
  NOR2_X1 U1339 ( .A1(n189), .A2(n281), .ZN(ab_11__10_) );
  NOR2_X1 U1340 ( .A1(n219), .A2(n281), .ZN(ab_11__0_) );
  NOR2_X1 U1341 ( .A1(n192), .A2(n286), .ZN(ab_10__9_) );
  NOR2_X1 U1342 ( .A1(n195), .A2(n286), .ZN(ab_10__8_) );
  NOR2_X1 U1343 ( .A1(n198), .A2(n286), .ZN(ab_10__7_) );
  NOR2_X1 U1344 ( .A1(n201), .A2(n286), .ZN(ab_10__6_) );
  NOR2_X1 U1345 ( .A1(n204), .A2(n286), .ZN(ab_10__5_) );
  NOR2_X1 U1346 ( .A1(n207), .A2(n286), .ZN(ab_10__4_) );
  NOR2_X1 U1347 ( .A1(n210), .A2(n286), .ZN(ab_10__3_) );
  NOR2_X1 U1348 ( .A1(A[10]), .A2(n127), .ZN(ab_10__31_) );
  NOR2_X1 U1349 ( .A1(n129), .A2(n285), .ZN(ab_10__30_) );
  NOR2_X1 U1350 ( .A1(n213), .A2(n285), .ZN(ab_10__2_) );
  NOR2_X1 U1351 ( .A1(n132), .A2(n285), .ZN(ab_10__29_) );
  NOR2_X1 U1352 ( .A1(n135), .A2(n285), .ZN(ab_10__28_) );
  NOR2_X1 U1353 ( .A1(n138), .A2(n285), .ZN(ab_10__27_) );
  NOR2_X1 U1354 ( .A1(n141), .A2(n285), .ZN(ab_10__26_) );
  NOR2_X1 U1355 ( .A1(n144), .A2(n285), .ZN(ab_10__25_) );
  NOR2_X1 U1356 ( .A1(n147), .A2(n285), .ZN(ab_10__24_) );
  NOR2_X1 U1357 ( .A1(n150), .A2(n285), .ZN(ab_10__23_) );
  NOR2_X1 U1358 ( .A1(n153), .A2(n285), .ZN(ab_10__22_) );
  NOR2_X1 U1359 ( .A1(n156), .A2(n285), .ZN(ab_10__21_) );
  NOR2_X1 U1360 ( .A1(n159), .A2(n285), .ZN(ab_10__20_) );
  NOR2_X1 U1361 ( .A1(n216), .A2(n284), .ZN(ab_10__1_) );
  NOR2_X1 U1362 ( .A1(n162), .A2(n284), .ZN(ab_10__19_) );
  NOR2_X1 U1363 ( .A1(n165), .A2(n284), .ZN(ab_10__18_) );
  NOR2_X1 U1364 ( .A1(n168), .A2(n284), .ZN(ab_10__17_) );
  NOR2_X1 U1365 ( .A1(n171), .A2(n284), .ZN(ab_10__16_) );
  NOR2_X1 U1366 ( .A1(n174), .A2(n284), .ZN(ab_10__15_) );
  NOR2_X1 U1367 ( .A1(n177), .A2(n284), .ZN(ab_10__14_) );
  NOR2_X1 U1368 ( .A1(n180), .A2(n284), .ZN(ab_10__13_) );
  NOR2_X1 U1369 ( .A1(n183), .A2(n284), .ZN(ab_10__12_) );
  NOR2_X1 U1370 ( .A1(n186), .A2(n284), .ZN(ab_10__11_) );
  NOR2_X1 U1371 ( .A1(n189), .A2(n284), .ZN(ab_10__10_) );
  NOR2_X1 U1372 ( .A1(n219), .A2(n284), .ZN(ab_10__0_) );
  NOR2_X1 U1373 ( .A1(n192), .A2(n316), .ZN(ab_0__9_) );
  NOR2_X1 U1374 ( .A1(n195), .A2(n316), .ZN(ab_0__8_) );
  NOR2_X1 U1375 ( .A1(n198), .A2(n316), .ZN(ab_0__7_) );
  NOR2_X1 U1376 ( .A1(n201), .A2(n316), .ZN(ab_0__6_) );
  NOR2_X1 U1377 ( .A1(n204), .A2(n316), .ZN(ab_0__5_) );
  NOR2_X1 U1378 ( .A1(n207), .A2(n316), .ZN(ab_0__4_) );
  NOR2_X1 U1379 ( .A1(n210), .A2(n316), .ZN(ab_0__3_) );
  NOR2_X1 U1380 ( .A1(A[0]), .A2(n127), .ZN(ab_0__31_) );
  NOR2_X1 U1381 ( .A1(n129), .A2(n315), .ZN(ab_0__30_) );
  NOR2_X1 U1382 ( .A1(n213), .A2(n315), .ZN(ab_0__2_) );
  NOR2_X1 U1383 ( .A1(n132), .A2(n315), .ZN(ab_0__29_) );
  NOR2_X1 U1384 ( .A1(n135), .A2(n315), .ZN(ab_0__28_) );
  NOR2_X1 U1385 ( .A1(n138), .A2(n315), .ZN(ab_0__27_) );
  NOR2_X1 U1386 ( .A1(n141), .A2(n315), .ZN(ab_0__26_) );
  NOR2_X1 U1387 ( .A1(n144), .A2(n315), .ZN(ab_0__25_) );
  NOR2_X1 U1388 ( .A1(n147), .A2(n315), .ZN(ab_0__24_) );
  NOR2_X1 U1389 ( .A1(n150), .A2(n315), .ZN(ab_0__23_) );
  NOR2_X1 U1390 ( .A1(n153), .A2(n315), .ZN(ab_0__22_) );
  NOR2_X1 U1391 ( .A1(n156), .A2(n315), .ZN(ab_0__21_) );
  NOR2_X1 U1392 ( .A1(n159), .A2(n315), .ZN(ab_0__20_) );
  NOR2_X1 U1393 ( .A1(n216), .A2(n314), .ZN(ab_0__1_) );
  NOR2_X1 U1394 ( .A1(n162), .A2(n314), .ZN(ab_0__19_) );
  NOR2_X1 U1395 ( .A1(n165), .A2(n314), .ZN(ab_0__18_) );
  NOR2_X1 U1396 ( .A1(n168), .A2(n314), .ZN(ab_0__17_) );
  NOR2_X1 U1397 ( .A1(n171), .A2(n314), .ZN(ab_0__16_) );
  NOR2_X1 U1398 ( .A1(n174), .A2(n314), .ZN(ab_0__15_) );
  NOR2_X1 U1399 ( .A1(n177), .A2(n314), .ZN(ab_0__14_) );
  NOR2_X1 U1400 ( .A1(n180), .A2(n314), .ZN(ab_0__13_) );
  NOR2_X1 U1401 ( .A1(n183), .A2(n314), .ZN(ab_0__12_) );
  NOR2_X1 U1402 ( .A1(n186), .A2(n314), .ZN(ab_0__11_) );
  NOR2_X1 U1403 ( .A1(n189), .A2(n314), .ZN(ab_0__10_) );
  NOR2_X1 U1404 ( .A1(n219), .A2(n314), .ZN(PRODUCT[0]) );
endmodule


module simpleMultiplier ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;


  simpleMultiplier_DW02_mult_0 mult_8 ( .A(a), .B(b), .TC(1'b1), .PRODUCT(
        result) );
endmodule


module register_N64 ( clk, reset, reg_in, reg_out );
  input [63:0] reg_in;
  output [63:0] reg_out;
  input clk, reset;
  wire   n83, n84, n85, n86, n87, n88, n89, n90, n91;

  SDFF_X1 reg_out_reg_63_ ( .D(1'b0), .SI(n85), .SE(reg_in[63]), .CK(clk), .Q(
        reg_out[63]) );
  SDFF_X1 reg_out_reg_62_ ( .D(1'b0), .SI(n85), .SE(reg_in[62]), .CK(clk), .Q(
        reg_out[62]) );
  SDFF_X1 reg_out_reg_61_ ( .D(1'b0), .SI(n85), .SE(reg_in[61]), .CK(clk), .Q(
        reg_out[61]) );
  SDFF_X1 reg_out_reg_60_ ( .D(1'b0), .SI(n85), .SE(reg_in[60]), .CK(clk), .Q(
        reg_out[60]) );
  SDFF_X1 reg_out_reg_59_ ( .D(1'b0), .SI(n85), .SE(reg_in[59]), .CK(clk), .Q(
        reg_out[59]) );
  SDFF_X1 reg_out_reg_58_ ( .D(1'b0), .SI(n85), .SE(reg_in[58]), .CK(clk), .Q(
        reg_out[58]) );
  SDFF_X1 reg_out_reg_57_ ( .D(1'b0), .SI(n85), .SE(reg_in[57]), .CK(clk), .Q(
        reg_out[57]) );
  SDFF_X1 reg_out_reg_56_ ( .D(1'b0), .SI(n85), .SE(reg_in[56]), .CK(clk), .Q(
        reg_out[56]) );
  SDFF_X1 reg_out_reg_55_ ( .D(1'b0), .SI(n85), .SE(reg_in[55]), .CK(clk), .Q(
        reg_out[55]) );
  SDFF_X1 reg_out_reg_54_ ( .D(1'b0), .SI(n85), .SE(reg_in[54]), .CK(clk), .Q(
        reg_out[54]) );
  SDFF_X1 reg_out_reg_53_ ( .D(1'b0), .SI(n85), .SE(reg_in[53]), .CK(clk), .Q(
        reg_out[53]) );
  SDFF_X1 reg_out_reg_52_ ( .D(1'b0), .SI(n84), .SE(reg_in[52]), .CK(clk), .Q(
        reg_out[52]) );
  SDFF_X1 reg_out_reg_51_ ( .D(1'b0), .SI(n84), .SE(reg_in[51]), .CK(clk), .Q(
        reg_out[51]) );
  SDFF_X1 reg_out_reg_50_ ( .D(1'b0), .SI(n84), .SE(reg_in[50]), .CK(clk), .Q(
        reg_out[50]) );
  SDFF_X1 reg_out_reg_49_ ( .D(1'b0), .SI(n84), .SE(reg_in[49]), .CK(clk), .Q(
        reg_out[49]) );
  SDFF_X1 reg_out_reg_48_ ( .D(1'b0), .SI(n84), .SE(reg_in[48]), .CK(clk), .Q(
        reg_out[48]) );
  SDFF_X1 reg_out_reg_47_ ( .D(1'b0), .SI(n84), .SE(reg_in[47]), .CK(clk), .Q(
        reg_out[47]) );
  SDFF_X1 reg_out_reg_46_ ( .D(1'b0), .SI(n84), .SE(reg_in[46]), .CK(clk), .Q(
        reg_out[46]) );
  SDFF_X1 reg_out_reg_45_ ( .D(1'b0), .SI(n84), .SE(reg_in[45]), .CK(clk), .Q(
        reg_out[45]) );
  SDFF_X1 reg_out_reg_44_ ( .D(1'b0), .SI(n84), .SE(reg_in[44]), .CK(clk), .Q(
        reg_out[44]) );
  SDFF_X1 reg_out_reg_43_ ( .D(1'b0), .SI(n84), .SE(reg_in[43]), .CK(clk), .Q(
        reg_out[43]) );
  SDFF_X1 reg_out_reg_42_ ( .D(1'b0), .SI(n84), .SE(reg_in[42]), .CK(clk), .Q(
        reg_out[42]) );
  SDFF_X1 reg_out_reg_41_ ( .D(1'b0), .SI(n83), .SE(reg_in[41]), .CK(clk), .Q(
        reg_out[41]) );
  SDFF_X1 reg_out_reg_40_ ( .D(1'b0), .SI(n83), .SE(reg_in[40]), .CK(clk), .Q(
        reg_out[40]) );
  SDFF_X1 reg_out_reg_39_ ( .D(1'b0), .SI(n83), .SE(reg_in[39]), .CK(clk), .Q(
        reg_out[39]) );
  SDFF_X1 reg_out_reg_38_ ( .D(1'b0), .SI(n83), .SE(reg_in[38]), .CK(clk), .Q(
        reg_out[38]) );
  SDFF_X1 reg_out_reg_37_ ( .D(1'b0), .SI(n83), .SE(reg_in[37]), .CK(clk), .Q(
        reg_out[37]) );
  SDFF_X1 reg_out_reg_36_ ( .D(1'b0), .SI(n83), .SE(reg_in[36]), .CK(clk), .Q(
        reg_out[36]) );
  SDFF_X1 reg_out_reg_35_ ( .D(1'b0), .SI(n83), .SE(reg_in[35]), .CK(clk), .Q(
        reg_out[35]) );
  SDFF_X1 reg_out_reg_34_ ( .D(1'b0), .SI(n83), .SE(reg_in[34]), .CK(clk), .Q(
        reg_out[34]) );
  SDFF_X1 reg_out_reg_33_ ( .D(1'b0), .SI(n83), .SE(reg_in[33]), .CK(clk), .Q(
        reg_out[33]) );
  SDFF_X1 reg_out_reg_32_ ( .D(1'b0), .SI(n83), .SE(reg_in[32]), .CK(clk), .Q(
        reg_out[32]) );
  SDFF_X1 reg_out_reg_31_ ( .D(1'b0), .SI(n83), .SE(reg_in[31]), .CK(clk), .Q(
        reg_out[31]) );
  SDFF_X1 reg_out_reg_30_ ( .D(1'b0), .SI(n87), .SE(reg_in[30]), .CK(clk), .Q(
        reg_out[30]) );
  SDFF_X1 reg_out_reg_29_ ( .D(1'b0), .SI(n87), .SE(reg_in[29]), .CK(clk), .Q(
        reg_out[29]) );
  SDFF_X1 reg_out_reg_28_ ( .D(1'b0), .SI(n87), .SE(reg_in[28]), .CK(clk), .Q(
        reg_out[28]) );
  SDFF_X1 reg_out_reg_27_ ( .D(1'b0), .SI(n87), .SE(reg_in[27]), .CK(clk), .Q(
        reg_out[27]) );
  SDFF_X1 reg_out_reg_26_ ( .D(1'b0), .SI(n87), .SE(reg_in[26]), .CK(clk), .Q(
        reg_out[26]) );
  SDFF_X1 reg_out_reg_25_ ( .D(1'b0), .SI(n87), .SE(reg_in[25]), .CK(clk), .Q(
        reg_out[25]) );
  SDFF_X1 reg_out_reg_24_ ( .D(1'b0), .SI(n87), .SE(reg_in[24]), .CK(clk), .Q(
        reg_out[24]) );
  SDFF_X1 reg_out_reg_23_ ( .D(1'b0), .SI(n87), .SE(reg_in[23]), .CK(clk), .Q(
        reg_out[23]) );
  SDFF_X1 reg_out_reg_22_ ( .D(1'b0), .SI(n87), .SE(reg_in[22]), .CK(clk), .Q(
        reg_out[22]) );
  SDFF_X1 reg_out_reg_21_ ( .D(1'b0), .SI(n87), .SE(reg_in[21]), .CK(clk), .Q(
        reg_out[21]) );
  SDFF_X1 reg_out_reg_20_ ( .D(1'b0), .SI(n87), .SE(reg_in[20]), .CK(clk), .Q(
        reg_out[20]) );
  SDFF_X1 reg_out_reg_19_ ( .D(1'b0), .SI(n86), .SE(reg_in[19]), .CK(clk), .Q(
        reg_out[19]) );
  SDFF_X1 reg_out_reg_18_ ( .D(1'b0), .SI(n86), .SE(reg_in[18]), .CK(clk), .Q(
        reg_out[18]) );
  SDFF_X1 reg_out_reg_17_ ( .D(1'b0), .SI(n86), .SE(reg_in[17]), .CK(clk), .Q(
        reg_out[17]) );
  SDFF_X1 reg_out_reg_16_ ( .D(1'b0), .SI(n86), .SE(reg_in[16]), .CK(clk), .Q(
        reg_out[16]) );
  SDFF_X1 reg_out_reg_15_ ( .D(1'b0), .SI(n86), .SE(reg_in[15]), .CK(clk), .Q(
        reg_out[15]) );
  SDFF_X1 reg_out_reg_14_ ( .D(1'b0), .SI(n86), .SE(reg_in[14]), .CK(clk), .Q(
        reg_out[14]) );
  SDFF_X1 reg_out_reg_13_ ( .D(1'b0), .SI(n86), .SE(reg_in[13]), .CK(clk), .Q(
        reg_out[13]) );
  SDFF_X1 reg_out_reg_12_ ( .D(1'b0), .SI(n86), .SE(reg_in[12]), .CK(clk), .Q(
        reg_out[12]) );
  SDFF_X1 reg_out_reg_11_ ( .D(1'b0), .SI(n86), .SE(reg_in[11]), .CK(clk), .Q(
        reg_out[11]) );
  SDFF_X1 reg_out_reg_10_ ( .D(1'b0), .SI(n86), .SE(reg_in[10]), .CK(clk), .Q(
        reg_out[10]) );
  SDFF_X1 reg_out_reg_9_ ( .D(1'b0), .SI(n86), .SE(reg_in[9]), .CK(clk), .Q(
        reg_out[9]) );
  SDFF_X1 reg_out_reg_8_ ( .D(1'b0), .SI(n88), .SE(reg_in[8]), .CK(clk), .Q(
        reg_out[8]) );
  SDFF_X1 reg_out_reg_7_ ( .D(1'b0), .SI(n88), .SE(reg_in[7]), .CK(clk), .Q(
        reg_out[7]) );
  SDFF_X1 reg_out_reg_6_ ( .D(1'b0), .SI(n88), .SE(reg_in[6]), .CK(clk), .Q(
        reg_out[6]) );
  SDFF_X1 reg_out_reg_5_ ( .D(1'b0), .SI(n88), .SE(reg_in[5]), .CK(clk), .Q(
        reg_out[5]) );
  SDFF_X1 reg_out_reg_4_ ( .D(1'b0), .SI(n88), .SE(reg_in[4]), .CK(clk), .Q(
        reg_out[4]) );
  SDFF_X1 reg_out_reg_3_ ( .D(1'b0), .SI(n88), .SE(reg_in[3]), .CK(clk), .Q(
        reg_out[3]) );
  SDFF_X1 reg_out_reg_2_ ( .D(1'b0), .SI(n88), .SE(reg_in[2]), .CK(clk), .Q(
        reg_out[2]) );
  SDFF_X1 reg_out_reg_1_ ( .D(1'b0), .SI(n88), .SE(reg_in[1]), .CK(clk), .Q(
        reg_out[1]) );
  SDFF_X1 reg_out_reg_0_ ( .D(1'b0), .SI(n88), .SE(reg_in[0]), .CK(clk), .Q(
        reg_out[0]) );
  BUF_X1 U67 ( .A(n89), .Z(n86) );
  BUF_X1 U68 ( .A(n89), .Z(n87) );
  BUF_X1 U69 ( .A(n90), .Z(n83) );
  BUF_X1 U70 ( .A(n90), .Z(n84) );
  BUF_X1 U71 ( .A(n90), .Z(n85) );
  BUF_X1 U72 ( .A(n89), .Z(n88) );
  INV_X1 U73 ( .A(reset), .ZN(n91) );
  BUF_X1 U74 ( .A(n91), .Z(n89) );
  BUF_X1 U75 ( .A(n91), .Z(n90) );
endmodule


module TopModule ( clk, a, b, reset, resetReg, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;
  input clk, reset, resetReg;

  wire   [31:0] mulA;
  wire   [31:0] mulB;
  wire   [63:0] mulResult;

  register_N32_2 R0 ( .clk(clk), .reset(resetReg), .reg_in(a), .reg_out(mulA)
         );
  register_N32_3 R1 ( .clk(clk), .reset(resetReg), .reg_in(b), .reg_out(mulB)
         );
  simpleMultiplier M0 ( .a(mulA), .b(mulB), .result(mulResult) );
  register_N64 R2 ( .clk(clk), .reset(resetReg), .reg_in(mulResult), .reg_out(
        result) );
endmodule

