
module register_N64_0 ( clk, reset, reg_in, reg_out );
  input [63:0] reg_in;
  output [63:0] reg_out;
  input clk, reset;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73;

  SDFF_X1 reg_out_reg_63_ ( .D(1'b0), .SI(n65), .SE(reg_in[63]), .CK(clk), .Q(
        reg_out[63]) );
  SDFF_X1 reg_out_reg_62_ ( .D(1'b0), .SI(n65), .SE(reg_in[62]), .CK(clk), .Q(
        reg_out[62]) );
  SDFF_X1 reg_out_reg_61_ ( .D(1'b0), .SI(n65), .SE(reg_in[61]), .CK(clk), .Q(
        reg_out[61]) );
  SDFF_X1 reg_out_reg_60_ ( .D(1'b0), .SI(n65), .SE(reg_in[60]), .CK(clk), .Q(
        reg_out[60]) );
  SDFF_X1 reg_out_reg_59_ ( .D(1'b0), .SI(n65), .SE(reg_in[59]), .CK(clk), .Q(
        reg_out[59]) );
  SDFF_X1 reg_out_reg_58_ ( .D(1'b0), .SI(n65), .SE(reg_in[58]), .CK(clk), .Q(
        reg_out[58]) );
  SDFF_X1 reg_out_reg_57_ ( .D(1'b0), .SI(n65), .SE(reg_in[57]), .CK(clk), .Q(
        reg_out[57]) );
  SDFF_X1 reg_out_reg_56_ ( .D(1'b0), .SI(n65), .SE(reg_in[56]), .CK(clk), .Q(
        reg_out[56]) );
  SDFF_X1 reg_out_reg_55_ ( .D(1'b0), .SI(n65), .SE(reg_in[55]), .CK(clk), .Q(
        reg_out[55]) );
  SDFF_X1 reg_out_reg_54_ ( .D(1'b0), .SI(n65), .SE(reg_in[54]), .CK(clk), .Q(
        reg_out[54]) );
  SDFF_X1 reg_out_reg_53_ ( .D(1'b0), .SI(n65), .SE(reg_in[53]), .CK(clk), .Q(
        reg_out[53]) );
  SDFF_X1 reg_out_reg_52_ ( .D(1'b0), .SI(n66), .SE(reg_in[52]), .CK(clk), .Q(
        reg_out[52]) );
  SDFF_X1 reg_out_reg_51_ ( .D(1'b0), .SI(n66), .SE(reg_in[51]), .CK(clk), .Q(
        reg_out[51]) );
  SDFF_X1 reg_out_reg_50_ ( .D(1'b0), .SI(n66), .SE(reg_in[50]), .CK(clk), .Q(
        reg_out[50]) );
  SDFF_X1 reg_out_reg_49_ ( .D(1'b0), .SI(n66), .SE(reg_in[49]), .CK(clk), .Q(
        reg_out[49]) );
  SDFF_X1 reg_out_reg_48_ ( .D(1'b0), .SI(n66), .SE(reg_in[48]), .CK(clk), .Q(
        reg_out[48]) );
  SDFF_X1 reg_out_reg_47_ ( .D(1'b0), .SI(n66), .SE(reg_in[47]), .CK(clk), .Q(
        reg_out[47]) );
  SDFF_X1 reg_out_reg_46_ ( .D(1'b0), .SI(n66), .SE(reg_in[46]), .CK(clk), .Q(
        reg_out[46]) );
  SDFF_X1 reg_out_reg_45_ ( .D(1'b0), .SI(n66), .SE(reg_in[45]), .CK(clk), .Q(
        reg_out[45]) );
  SDFF_X1 reg_out_reg_44_ ( .D(1'b0), .SI(n66), .SE(reg_in[44]), .CK(clk), .Q(
        reg_out[44]) );
  SDFF_X1 reg_out_reg_43_ ( .D(1'b0), .SI(n66), .SE(reg_in[43]), .CK(clk), .Q(
        reg_out[43]) );
  SDFF_X1 reg_out_reg_42_ ( .D(1'b0), .SI(n66), .SE(reg_in[42]), .CK(clk), .Q(
        reg_out[42]) );
  SDFF_X1 reg_out_reg_41_ ( .D(1'b0), .SI(n67), .SE(reg_in[41]), .CK(clk), .Q(
        reg_out[41]) );
  SDFF_X1 reg_out_reg_40_ ( .D(1'b0), .SI(n67), .SE(reg_in[40]), .CK(clk), .Q(
        reg_out[40]) );
  SDFF_X1 reg_out_reg_39_ ( .D(1'b0), .SI(n67), .SE(reg_in[39]), .CK(clk), .Q(
        reg_out[39]) );
  SDFF_X1 reg_out_reg_38_ ( .D(1'b0), .SI(n67), .SE(reg_in[38]), .CK(clk), .Q(
        reg_out[38]) );
  SDFF_X1 reg_out_reg_37_ ( .D(1'b0), .SI(n67), .SE(reg_in[37]), .CK(clk), .Q(
        reg_out[37]) );
  SDFF_X1 reg_out_reg_36_ ( .D(1'b0), .SI(n67), .SE(reg_in[36]), .CK(clk), .Q(
        reg_out[36]) );
  SDFF_X1 reg_out_reg_35_ ( .D(1'b0), .SI(n67), .SE(reg_in[35]), .CK(clk), .Q(
        reg_out[35]) );
  SDFF_X1 reg_out_reg_34_ ( .D(1'b0), .SI(n67), .SE(reg_in[34]), .CK(clk), .Q(
        reg_out[34]) );
  SDFF_X1 reg_out_reg_33_ ( .D(1'b0), .SI(n67), .SE(reg_in[33]), .CK(clk), .Q(
        reg_out[33]) );
  SDFF_X1 reg_out_reg_32_ ( .D(1'b0), .SI(n67), .SE(reg_in[32]), .CK(clk), .Q(
        reg_out[32]) );
  SDFF_X1 reg_out_reg_31_ ( .D(1'b0), .SI(n67), .SE(reg_in[31]), .CK(clk), .Q(
        reg_out[31]) );
  SDFF_X1 reg_out_reg_30_ ( .D(1'b0), .SI(n68), .SE(reg_in[30]), .CK(clk), .Q(
        reg_out[30]) );
  SDFF_X1 reg_out_reg_29_ ( .D(1'b0), .SI(n68), .SE(reg_in[29]), .CK(clk), .Q(
        reg_out[29]) );
  SDFF_X1 reg_out_reg_28_ ( .D(1'b0), .SI(n68), .SE(reg_in[28]), .CK(clk), .Q(
        reg_out[28]) );
  SDFF_X1 reg_out_reg_27_ ( .D(1'b0), .SI(n68), .SE(reg_in[27]), .CK(clk), .Q(
        reg_out[27]) );
  SDFF_X1 reg_out_reg_26_ ( .D(1'b0), .SI(n68), .SE(reg_in[26]), .CK(clk), .Q(
        reg_out[26]) );
  SDFF_X1 reg_out_reg_25_ ( .D(1'b0), .SI(n68), .SE(reg_in[25]), .CK(clk), .Q(
        reg_out[25]) );
  SDFF_X1 reg_out_reg_24_ ( .D(1'b0), .SI(n68), .SE(reg_in[24]), .CK(clk), .Q(
        reg_out[24]) );
  SDFF_X1 reg_out_reg_23_ ( .D(1'b0), .SI(n68), .SE(reg_in[23]), .CK(clk), .Q(
        reg_out[23]) );
  SDFF_X1 reg_out_reg_22_ ( .D(1'b0), .SI(n68), .SE(reg_in[22]), .CK(clk), .Q(
        reg_out[22]) );
  SDFF_X1 reg_out_reg_21_ ( .D(1'b0), .SI(n68), .SE(reg_in[21]), .CK(clk), .Q(
        reg_out[21]) );
  SDFF_X1 reg_out_reg_20_ ( .D(1'b0), .SI(n68), .SE(reg_in[20]), .CK(clk), .Q(
        reg_out[20]) );
  SDFF_X1 reg_out_reg_19_ ( .D(1'b0), .SI(n69), .SE(reg_in[19]), .CK(clk), .Q(
        reg_out[19]) );
  SDFF_X1 reg_out_reg_18_ ( .D(1'b0), .SI(n69), .SE(reg_in[18]), .CK(clk), .Q(
        reg_out[18]) );
  SDFF_X1 reg_out_reg_17_ ( .D(1'b0), .SI(n69), .SE(reg_in[17]), .CK(clk), .Q(
        reg_out[17]) );
  SDFF_X1 reg_out_reg_16_ ( .D(1'b0), .SI(n69), .SE(reg_in[16]), .CK(clk), .Q(
        reg_out[16]) );
  SDFF_X1 reg_out_reg_15_ ( .D(1'b0), .SI(n69), .SE(reg_in[15]), .CK(clk), .Q(
        reg_out[15]) );
  SDFF_X1 reg_out_reg_14_ ( .D(1'b0), .SI(n69), .SE(reg_in[14]), .CK(clk), .Q(
        reg_out[14]) );
  SDFF_X1 reg_out_reg_13_ ( .D(1'b0), .SI(n69), .SE(reg_in[13]), .CK(clk), .Q(
        reg_out[13]) );
  SDFF_X1 reg_out_reg_12_ ( .D(1'b0), .SI(n69), .SE(reg_in[12]), .CK(clk), .Q(
        reg_out[12]) );
  SDFF_X1 reg_out_reg_11_ ( .D(1'b0), .SI(n69), .SE(reg_in[11]), .CK(clk), .Q(
        reg_out[11]) );
  SDFF_X1 reg_out_reg_10_ ( .D(1'b0), .SI(n69), .SE(reg_in[10]), .CK(clk), .Q(
        reg_out[10]) );
  SDFF_X1 reg_out_reg_9_ ( .D(1'b0), .SI(n69), .SE(reg_in[9]), .CK(clk), .Q(
        reg_out[9]) );
  SDFF_X1 reg_out_reg_8_ ( .D(1'b0), .SI(n70), .SE(reg_in[8]), .CK(clk), .Q(
        reg_out[8]) );
  SDFF_X1 reg_out_reg_7_ ( .D(1'b0), .SI(n70), .SE(reg_in[7]), .CK(clk), .Q(
        reg_out[7]) );
  SDFF_X1 reg_out_reg_6_ ( .D(1'b0), .SI(n70), .SE(reg_in[6]), .CK(clk), .Q(
        reg_out[6]) );
  SDFF_X1 reg_out_reg_5_ ( .D(1'b0), .SI(n70), .SE(reg_in[5]), .CK(clk), .Q(
        reg_out[5]) );
  SDFF_X1 reg_out_reg_4_ ( .D(1'b0), .SI(n70), .SE(reg_in[4]), .CK(clk), .Q(
        reg_out[4]) );
  SDFF_X1 reg_out_reg_3_ ( .D(1'b0), .SI(n70), .SE(reg_in[3]), .CK(clk), .Q(
        reg_out[3]) );
  SDFF_X1 reg_out_reg_2_ ( .D(1'b0), .SI(n70), .SE(reg_in[2]), .CK(clk), .Q(
        reg_out[2]) );
  SDFF_X1 reg_out_reg_1_ ( .D(1'b0), .SI(n70), .SE(reg_in[1]), .CK(clk), .Q(
        reg_out[1]) );
  SDFF_X1 reg_out_reg_0_ ( .D(1'b0), .SI(n70), .SE(reg_in[0]), .CK(clk), .Q(
        reg_out[0]) );
  BUF_X1 U67 ( .A(n71), .Z(n69) );
  BUF_X1 U68 ( .A(n71), .Z(n68) );
  BUF_X1 U69 ( .A(n72), .Z(n66) );
  BUF_X1 U70 ( .A(n72), .Z(n65) );
  BUF_X1 U71 ( .A(n71), .Z(n70) );
  INV_X1 U72 ( .A(reset), .ZN(n73) );
  BUF_X1 U73 ( .A(n72), .Z(n67) );
  BUF_X1 U74 ( .A(n73), .Z(n71) );
  BUF_X1 U75 ( .A(n73), .Z(n72) );
endmodule


module carryLookAheadAdder64bit ( a, b, cin, result, cout );
  input [63:0] a;
  input [63:0] b;
  output [63:0] result;
  input cin;
  output cout;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n132, n134, n136, n138, n140, n141, n143, n145,
         n146, n147, n149, n151, n152, n154, n156, n158, n160, n162, n164,
         n165, n167, n168, n170, n171, n172, n174, n175, n177, n178, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n131, n133, n135, n137, n139, n142,
         n144, n148, n150, n153, n155, n157, n159, n161, n163, n166, n169,
         n173, n176, n179, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273;

  XOR2_X1 U130 ( .A(n265), .B(n67), .Z(result[8]) );
  XOR2_X1 U131 ( .A(n68), .B(n266), .Z(result[7]) );
  XOR2_X1 U132 ( .A(n267), .B(n69), .Z(result[6]) );
  XOR2_X1 U134 ( .A(n44), .B(n72), .Z(result[62]) );
  XOR2_X1 U135 ( .A(n73), .B(n231), .Z(result[61]) );
  XOR2_X1 U136 ( .A(n39), .B(n74), .Z(result[60]) );
  XOR2_X1 U137 ( .A(n75), .B(n268), .Z(result[5]) );
  XOR2_X1 U138 ( .A(n76), .B(n232), .Z(result[59]) );
  XOR2_X1 U139 ( .A(n22), .B(n77), .Z(result[58]) );
  XOR2_X1 U140 ( .A(n78), .B(n233), .Z(result[57]) );
  XOR2_X1 U141 ( .A(n53), .B(n79), .Z(result[56]) );
  XOR2_X1 U142 ( .A(n234), .B(n80), .Z(result[55]) );
  XOR2_X1 U143 ( .A(n135), .B(n81), .Z(result[54]) );
  XOR2_X1 U144 ( .A(n82), .B(n235), .Z(result[53]) );
  XOR2_X1 U145 ( .A(n236), .B(n83), .Z(result[52]) );
  XOR2_X1 U146 ( .A(n84), .B(n17), .Z(result[51]) );
  XOR2_X1 U147 ( .A(n237), .B(n85), .Z(result[50]) );
  XOR2_X1 U148 ( .A(n269), .B(n86), .Z(result[4]) );
  XOR2_X1 U149 ( .A(n87), .B(n16), .Z(result[49]) );
  XOR2_X1 U150 ( .A(n238), .B(n88), .Z(result[48]) );
  XOR2_X1 U151 ( .A(n89), .B(n64), .Z(result[47]) );
  XOR2_X1 U152 ( .A(n240), .B(n90), .Z(result[46]) );
  XOR2_X1 U153 ( .A(n91), .B(n19), .Z(result[45]) );
  XOR2_X1 U154 ( .A(n241), .B(n92), .Z(result[44]) );
  XOR2_X1 U155 ( .A(n93), .B(n18), .Z(result[43]) );
  XOR2_X1 U156 ( .A(n242), .B(n94), .Z(result[42]) );
  XOR2_X1 U157 ( .A(n95), .B(n243), .Z(result[41]) );
  XOR2_X1 U158 ( .A(n57), .B(n96), .Z(result[40]) );
  XOR2_X1 U159 ( .A(n97), .B(n63), .Z(result[3]) );
  XOR2_X1 U160 ( .A(n98), .B(n244), .Z(result[39]) );
  XOR2_X1 U161 ( .A(n7), .B(n99), .Z(result[38]) );
  XOR2_X1 U162 ( .A(n100), .B(n245), .Z(result[37]) );
  XOR2_X1 U163 ( .A(n49), .B(n101), .Z(result[36]) );
  XOR2_X1 U164 ( .A(n102), .B(n246), .Z(result[35]) );
  XOR2_X1 U165 ( .A(n13), .B(n103), .Z(result[34]) );
  XOR2_X1 U166 ( .A(n104), .B(n247), .Z(result[33]) );
  XOR2_X1 U167 ( .A(n11), .B(n105), .Z(result[32]) );
  XOR2_X1 U168 ( .A(n106), .B(n248), .Z(result[31]) );
  XOR2_X1 U169 ( .A(n6), .B(n107), .Z(result[30]) );
  XOR2_X1 U170 ( .A(n108), .B(n229), .Z(result[2]) );
  XOR2_X1 U171 ( .A(n109), .B(n249), .Z(result[29]) );
  XOR2_X1 U172 ( .A(n43), .B(n110), .Z(result[28]) );
  XOR2_X1 U173 ( .A(n111), .B(n20), .Z(result[27]) );
  XOR2_X1 U174 ( .A(n251), .B(n112), .Z(result[26]) );
  XOR2_X1 U175 ( .A(n113), .B(n252), .Z(result[25]) );
  XOR2_X1 U176 ( .A(n14), .B(n114), .Z(result[24]) );
  XOR2_X1 U177 ( .A(n115), .B(n253), .Z(result[23]) );
  XOR2_X1 U178 ( .A(n254), .B(n116), .Z(result[22]) );
  XOR2_X1 U179 ( .A(n117), .B(n255), .Z(result[21]) );
  XOR2_X1 U180 ( .A(n12), .B(n118), .Z(result[20]) );
  XOR2_X1 U181 ( .A(n119), .B(n272), .Z(result[1]) );
  XOR2_X1 U182 ( .A(n120), .B(n256), .Z(result[19]) );
  XOR2_X1 U183 ( .A(n257), .B(n121), .Z(result[18]) );
  XOR2_X1 U184 ( .A(n122), .B(n21), .Z(result[17]) );
  XOR2_X1 U185 ( .A(n258), .B(n123), .Z(result[16]) );
  XOR2_X1 U186 ( .A(n124), .B(n61), .Z(result[15]) );
  XOR2_X1 U187 ( .A(n15), .B(n125), .Z(result[14]) );
  XOR2_X1 U188 ( .A(n126), .B(n260), .Z(result[13]) );
  XOR2_X1 U189 ( .A(n261), .B(n127), .Z(result[12]) );
  XOR2_X1 U190 ( .A(n128), .B(n262), .Z(result[11]) );
  XOR2_X1 U191 ( .A(n263), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(cin), .B(n9), .Z(result[0]) );
  XOR2_X1 U193 ( .A(n273), .B(b[63]), .Z(n70) );
  XOR2_X1 U194 ( .A(a[62]), .B(b[62]), .Z(n72) );
  XOR2_X1 U196 ( .A(a[60]), .B(b[60]), .Z(n74) );
  XOR2_X1 U198 ( .A(a[58]), .B(b[58]), .Z(n77) );
  XOR2_X1 U200 ( .A(a[56]), .B(b[56]), .Z(n79) );
  XOR2_X1 U202 ( .A(a[54]), .B(b[54]), .Z(n81) );
  XOR2_X1 U204 ( .A(a[52]), .B(b[52]), .Z(n83) );
  XOR2_X1 U205 ( .A(a[51]), .B(b[51]), .Z(n84) );
  XOR2_X1 U207 ( .A(a[49]), .B(b[49]), .Z(n87) );
  XOR2_X1 U209 ( .A(a[47]), .B(b[47]), .Z(n89) );
  XOR2_X1 U210 ( .A(a[46]), .B(b[46]), .Z(n90) );
  XOR2_X1 U211 ( .A(a[45]), .B(b[45]), .Z(n91) );
  XOR2_X1 U213 ( .A(a[43]), .B(b[43]), .Z(n93) );
  XOR2_X1 U215 ( .A(a[41]), .B(b[41]), .Z(n95) );
  XOR2_X1 U216 ( .A(a[40]), .B(b[40]), .Z(n96) );
  XOR2_X1 U218 ( .A(a[38]), .B(b[38]), .Z(n99) );
  XOR2_X1 U220 ( .A(a[36]), .B(b[36]), .Z(n101) );
  XOR2_X1 U222 ( .A(a[34]), .B(b[34]), .Z(n103) );
  XOR2_X1 U223 ( .A(a[33]), .B(b[33]), .Z(n104) );
  XOR2_X1 U224 ( .A(a[32]), .B(b[32]), .Z(n105) );
  XOR2_X1 U226 ( .A(a[30]), .B(b[30]), .Z(n107) );
  XOR2_X1 U228 ( .A(a[28]), .B(b[28]), .Z(n110) );
  XOR2_X1 U229 ( .A(a[27]), .B(b[27]), .Z(n111) );
  XOR2_X1 U231 ( .A(a[25]), .B(b[25]), .Z(n113) );
  XOR2_X1 U232 ( .A(a[24]), .B(b[24]), .Z(n114) );
  XOR2_X1 U233 ( .A(a[23]), .B(b[23]), .Z(n115) );
  XOR2_X1 U234 ( .A(a[22]), .B(b[22]), .Z(n116) );
  XOR2_X1 U235 ( .A(a[21]), .B(b[21]), .Z(n117) );
  XOR2_X1 U236 ( .A(a[20]), .B(b[20]), .Z(n118) );
  XOR2_X1 U238 ( .A(a[18]), .B(b[18]), .Z(n121) );
  XOR2_X1 U239 ( .A(a[17]), .B(b[17]), .Z(n122) );
  XOR2_X1 U240 ( .A(a[16]), .B(b[16]), .Z(n123) );
  XOR2_X1 U241 ( .A(a[15]), .B(b[15]), .Z(n124) );
  XOR2_X1 U242 ( .A(a[14]), .B(b[14]), .Z(n125) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n126) );
  XOR2_X1 U244 ( .A(a[12]), .B(b[12]), .Z(n127) );
  XOR2_X1 U245 ( .A(a[11]), .B(b[11]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U247 ( .A(a[9]), .B(b[9]), .Z(n65) );
  XOR2_X1 U248 ( .A(a[8]), .B(b[8]), .Z(n67) );
  XOR2_X1 U249 ( .A(a[7]), .B(b[7]), .Z(n68) );
  XOR2_X1 U250 ( .A(a[6]), .B(b[6]), .Z(n69) );
  XOR2_X1 U251 ( .A(a[5]), .B(b[5]), .Z(n75) );
  XOR2_X1 U252 ( .A(a[4]), .B(b[4]), .Z(n86) );
  XOR2_X1 U253 ( .A(a[3]), .B(b[3]), .Z(n97) );
  XOR2_X1 U254 ( .A(a[2]), .B(b[2]), .Z(n108) );
  XOR2_X1 U255 ( .A(b[1]), .B(a[1]), .Z(n119) );
  XOR2_X1 U256 ( .A(b[0]), .B(a[0]), .Z(n130) );
  INV_X1 U1 ( .A(n73), .ZN(n48) );
  INV_X1 U2 ( .A(a[61]), .ZN(n47) );
  INV_X1 U3 ( .A(n76), .ZN(n155) );
  INV_X1 U4 ( .A(a[59]), .ZN(n153) );
  INV_X1 U5 ( .A(a[57]), .ZN(n214) );
  INV_X1 U6 ( .A(n78), .ZN(n215) );
  INV_X1 U7 ( .A(a[55]), .ZN(n55) );
  INV_X1 U8 ( .A(n80), .ZN(n56) );
  INV_X1 U9 ( .A(n82), .ZN(n176) );
  INV_X1 U10 ( .A(a[53]), .ZN(n173) );
  INV_X1 U11 ( .A(a[50]), .ZN(n33) );
  INV_X1 U12 ( .A(n85), .ZN(n34) );
  INV_X1 U13 ( .A(a[48]), .ZN(n161) );
  INV_X1 U14 ( .A(n88), .ZN(n163) );
  INV_X1 U15 ( .A(a[44]), .ZN(n25) );
  INV_X1 U16 ( .A(n92), .ZN(n26) );
  INV_X1 U17 ( .A(a[42]), .ZN(n193) );
  INV_X1 U18 ( .A(n94), .ZN(n194) );
  INV_X1 U19 ( .A(a[39]), .ZN(n59) );
  INV_X1 U20 ( .A(n98), .ZN(n60) );
  INV_X1 U21 ( .A(a[37]), .ZN(n198) );
  INV_X1 U22 ( .A(n100), .ZN(n199) );
  INV_X1 U23 ( .A(a[35]), .ZN(n51) );
  INV_X1 U24 ( .A(n102), .ZN(n52) );
  INV_X1 U25 ( .A(a[31]), .ZN(n29) );
  INV_X1 U26 ( .A(n106), .ZN(n30) );
  INV_X1 U27 ( .A(a[29]), .ZN(n142) );
  INV_X1 U28 ( .A(n109), .ZN(n144) );
  INV_X1 U29 ( .A(a[26]), .ZN(n202) );
  INV_X1 U30 ( .A(n112), .ZN(n203) );
  INV_X1 U31 ( .A(a[19]), .ZN(n210) );
  INV_X1 U32 ( .A(b[19]), .ZN(n209) );
  INV_X1 U33 ( .A(n120), .ZN(n211) );
  INV_X1 U34 ( .A(a[16]), .ZN(n206) );
  CLKBUF_X1 U35 ( .A(n134), .Z(n1) );
  CLKBUF_X1 U36 ( .A(n154), .Z(n2) );
  AOI22_X1 U37 ( .A1(b[58]), .A2(a[58]), .B1(n212), .B2(n77), .ZN(n134) );
  CLKBUF_X1 U38 ( .A(n138), .Z(n3) );
  CLKBUF_X1 U39 ( .A(n136), .Z(n4) );
  CLKBUF_X1 U40 ( .A(n143), .Z(n5) );
  CLKBUF_X1 U41 ( .A(n137), .Z(n6) );
  CLKBUF_X1 U42 ( .A(n196), .Z(n7) );
  AOI22_X1 U43 ( .A1(b[60]), .A2(a[60]), .B1(n148), .B2(n74), .ZN(n8) );
  CLKBUF_X1 U44 ( .A(n130), .Z(n9) );
  AOI22_X1 U45 ( .A1(b[8]), .A2(a[8]), .B1(n265), .B2(n67), .ZN(n10) );
  CLKBUF_X1 U46 ( .A(n27), .Z(n11) );
  CLKBUF_X1 U47 ( .A(n208), .Z(n12) );
  CLKBUF_X1 U48 ( .A(n225), .Z(n13) );
  CLKBUF_X1 U49 ( .A(n221), .Z(n14) );
  CLKBUF_X1 U50 ( .A(n217), .Z(n15) );
  CLKBUF_X1 U51 ( .A(n157), .Z(n16) );
  CLKBUF_X1 U52 ( .A(n31), .Z(n17) );
  CLKBUF_X1 U53 ( .A(n179), .Z(n18) );
  CLKBUF_X1 U54 ( .A(n23), .Z(n19) );
  CLKBUF_X1 U55 ( .A(n200), .Z(n20) );
  CLKBUF_X1 U56 ( .A(n204), .Z(n21) );
  CLKBUF_X1 U57 ( .A(n212), .Z(n22) );
  INV_X1 U58 ( .A(b[50]), .ZN(n32) );
  INV_X1 U59 ( .A(b[55]), .ZN(n54) );
  INV_X1 U60 ( .A(b[44]), .ZN(n24) );
  INV_X1 U61 ( .A(b[48]), .ZN(n159) );
  INV_X1 U62 ( .A(b[26]), .ZN(n201) );
  INV_X1 U63 ( .A(b[42]), .ZN(n192) );
  INV_X1 U64 ( .A(n70), .ZN(n62) );
  INV_X1 U65 ( .A(b[16]), .ZN(n205) );
  XOR2_X2 U66 ( .A(a[19]), .B(b[19]), .Z(n120) );
  INV_X1 U67 ( .A(b[29]), .ZN(n139) );
  XOR2_X2 U68 ( .A(a[29]), .B(b[29]), .Z(n109) );
  INV_X1 U69 ( .A(b[31]), .ZN(n28) );
  XOR2_X2 U70 ( .A(a[31]), .B(b[31]), .Z(n106) );
  INV_X1 U71 ( .A(b[35]), .ZN(n50) );
  XOR2_X2 U72 ( .A(a[35]), .B(b[35]), .Z(n102) );
  INV_X1 U73 ( .A(b[37]), .ZN(n197) );
  XOR2_X2 U74 ( .A(a[37]), .B(b[37]), .Z(n100) );
  INV_X1 U75 ( .A(b[39]), .ZN(n58) );
  XOR2_X2 U76 ( .A(a[39]), .B(b[39]), .Z(n98) );
  INV_X1 U77 ( .A(b[53]), .ZN(n169) );
  XOR2_X2 U78 ( .A(a[53]), .B(b[53]), .Z(n82) );
  INV_X1 U79 ( .A(b[57]), .ZN(n213) );
  XOR2_X2 U80 ( .A(a[57]), .B(b[57]), .Z(n78) );
  INV_X1 U81 ( .A(b[59]), .ZN(n150) );
  XOR2_X2 U82 ( .A(a[59]), .B(b[59]), .Z(n76) );
  INV_X1 U83 ( .A(b[61]), .ZN(n46) );
  XOR2_X2 U84 ( .A(a[61]), .B(b[61]), .Z(n73) );
  XOR2_X2 U85 ( .A(a[50]), .B(b[50]), .Z(n85) );
  XOR2_X2 U86 ( .A(a[55]), .B(b[55]), .Z(n80) );
  XOR2_X2 U87 ( .A(a[44]), .B(b[44]), .Z(n92) );
  XOR2_X2 U88 ( .A(a[48]), .B(b[48]), .Z(n88) );
  XOR2_X2 U89 ( .A(a[26]), .B(b[26]), .Z(n112) );
  XOR2_X2 U90 ( .A(a[42]), .B(b[42]), .Z(n94) );
  OAI22_X1 U91 ( .A1(n24), .A2(n25), .B1(n149), .B2(n26), .ZN(n23) );
  OAI22_X1 U92 ( .A1(n28), .A2(n29), .B1(n162), .B2(n30), .ZN(n27) );
  OAI22_X1 U93 ( .A1(n32), .A2(n33), .B1(n143), .B2(n34), .ZN(n31) );
  AOI22_X1 U94 ( .A1(b[52]), .A2(a[52]), .B1(n236), .B2(n83), .ZN(n35) );
  AOI22_X1 U95 ( .A1(b[41]), .A2(a[41]), .B1(n243), .B2(n95), .ZN(n36) );
  AOI22_X1 U96 ( .A1(b[22]), .A2(a[22]), .B1(n254), .B2(n116), .ZN(n37) );
  AOI22_X1 U97 ( .A1(b[25]), .A2(a[25]), .B1(n252), .B2(n113), .ZN(n38) );
  OAI22_X1 U98 ( .A1(n150), .A2(n153), .B1(n134), .B2(n155), .ZN(n39) );
  AOI22_X1 U99 ( .A1(b[52]), .A2(a[52]), .B1(n236), .B2(n83), .ZN(n140) );
  AOI22_X1 U100 ( .A1(b[18]), .A2(a[18]), .B1(n257), .B2(n121), .ZN(n40) );
  AOI22_X1 U101 ( .A1(b[12]), .A2(a[12]), .B1(n261), .B2(n127), .ZN(n41) );
  AOI22_X1 U102 ( .A1(b[60]), .A2(a[60]), .B1(n39), .B2(n74), .ZN(n42) );
  CLKBUF_X1 U103 ( .A(n250), .Z(n43) );
  OAI22_X1 U104 ( .A1(n46), .A2(n47), .B1(n42), .B2(n48), .ZN(n44) );
  OAI22_X1 U105 ( .A1(n46), .A2(n47), .B1(n8), .B2(n48), .ZN(n45) );
  OAI22_X1 U106 ( .A1(n50), .A2(n51), .B1(n158), .B2(n52), .ZN(n49) );
  OAI22_X1 U107 ( .A1(n54), .A2(n55), .B1(n138), .B2(n56), .ZN(n53) );
  OAI22_X1 U108 ( .A1(n58), .A2(n59), .B1(n154), .B2(n60), .ZN(n57) );
  INV_X1 U109 ( .A(n123), .ZN(n207) );
  CLKBUF_X1 U110 ( .A(n259), .Z(n61) );
  XNOR2_X1 U111 ( .A(n71), .B(n62), .ZN(result[63]) );
  CLKBUF_X1 U112 ( .A(n270), .Z(n63) );
  CLKBUF_X1 U113 ( .A(n239), .Z(n64) );
  AOI22_X1 U114 ( .A1(b[28]), .A2(a[28]), .B1(n43), .B2(n110), .ZN(n131) );
  AOI22_X1 U115 ( .A1(b[15]), .A2(a[15]), .B1(n61), .B2(n124), .ZN(n133) );
  OAI22_X1 U116 ( .A1(n169), .A2(n173), .B1(n35), .B2(n176), .ZN(n135) );
  OAI22_X1 U117 ( .A1(n139), .A2(n142), .B1(n164), .B2(n144), .ZN(n137) );
  OAI22_X1 U118 ( .A1(n150), .A2(n153), .B1(n134), .B2(n155), .ZN(n148) );
  OAI22_X1 U119 ( .A1(n159), .A2(n161), .B1(n145), .B2(n163), .ZN(n157) );
  OAI22_X1 U120 ( .A1(n169), .A2(n173), .B1(n140), .B2(n176), .ZN(n166) );
  OAI22_X1 U121 ( .A1(n192), .A2(n193), .B1(n151), .B2(n194), .ZN(n179) );
  AOI22_X1 U122 ( .A1(b[47]), .A2(a[47]), .B1(n64), .B2(n89), .ZN(n195) );
  OAI22_X1 U123 ( .A1(n197), .A2(n198), .B1(n156), .B2(n199), .ZN(n196) );
  OAI22_X1 U124 ( .A1(n201), .A2(n202), .B1(n167), .B2(n203), .ZN(n200) );
  OAI22_X1 U125 ( .A1(n205), .A2(n206), .B1(n177), .B2(n207), .ZN(n204) );
  OAI22_X1 U126 ( .A1(n209), .A2(n210), .B1(n174), .B2(n211), .ZN(n208) );
  OAI22_X1 U127 ( .A1(n213), .A2(n214), .B1(n136), .B2(n215), .ZN(n212) );
  INV_X1 U128 ( .A(b[63]), .ZN(n230) );
  INV_X1 U129 ( .A(a[23]), .ZN(n223) );
  INV_X1 U133 ( .A(b[23]), .ZN(n222) );
  INV_X1 U195 ( .A(n115), .ZN(n224) );
  INV_X1 U197 ( .A(a[33]), .ZN(n227) );
  INV_X1 U199 ( .A(b[33]), .ZN(n226) );
  INV_X1 U201 ( .A(n104), .ZN(n228) );
  INV_X1 U203 ( .A(a[13]), .ZN(n219) );
  INV_X1 U206 ( .A(b[13]), .ZN(n218) );
  INV_X1 U208 ( .A(a[63]), .ZN(n273) );
  AOI22_X1 U212 ( .A1(b[18]), .A2(a[18]), .B1(n257), .B2(n121), .ZN(n174) );
  AOI22_X1 U214 ( .A1(b[62]), .A2(a[62]), .B1(n44), .B2(n72), .ZN(n216) );
  INV_X1 U217 ( .A(n126), .ZN(n220) );
  OAI22_X1 U219 ( .A1(n218), .A2(n219), .B1(n180), .B2(n220), .ZN(n217) );
  AOI22_X1 U221 ( .A1(b[3]), .A2(a[3]), .B1(n270), .B2(n97), .ZN(n188) );
  OAI22_X1 U225 ( .A1(n222), .A2(n223), .B1(n170), .B2(n224), .ZN(n221) );
  OAI22_X1 U227 ( .A1(n226), .A2(n227), .B1(n160), .B2(n228), .ZN(n225) );
  CLKBUF_X1 U230 ( .A(n271), .Z(n229) );
  AOI22_X1 U237 ( .A1(b[1]), .A2(a[1]), .B1(n119), .B2(n272), .ZN(n190) );
  AOI22_X1 U257 ( .A1(b[2]), .A2(a[2]), .B1(n271), .B2(n108), .ZN(n189) );
  AOI22_X1 U258 ( .A1(b[28]), .A2(a[28]), .B1(n250), .B2(n110), .ZN(n164) );
  AOI22_X1 U259 ( .A1(b[43]), .A2(a[43]), .B1(n179), .B2(n93), .ZN(n149) );
  AOI22_X1 U260 ( .A1(b[4]), .A2(a[4]), .B1(n269), .B2(n86), .ZN(n187) );
  INV_X1 U261 ( .A(n188), .ZN(n269) );
  AOI22_X1 U262 ( .A1(b[38]), .A2(a[38]), .B1(n196), .B2(n99), .ZN(n154) );
  AOI22_X1 U263 ( .A1(b[27]), .A2(a[27]), .B1(n200), .B2(n111), .ZN(n165) );
  AOI22_X1 U264 ( .A1(b[17]), .A2(a[17]), .B1(n204), .B2(n122), .ZN(n175) );
  INV_X1 U265 ( .A(n190), .ZN(n271) );
  INV_X1 U266 ( .A(n189), .ZN(n270) );
  AOI22_X1 U267 ( .A1(b[49]), .A2(a[49]), .B1(n157), .B2(n87), .ZN(n143) );
  AOI22_X1 U268 ( .A1(b[7]), .A2(a[7]), .B1(n266), .B2(n68), .ZN(n184) );
  INV_X1 U269 ( .A(n132), .ZN(n231) );
  AOI22_X1 U270 ( .A1(b[47]), .A2(a[47]), .B1(n239), .B2(n89), .ZN(n145) );
  INV_X1 U271 ( .A(n160), .ZN(n247) );
  INV_X1 U272 ( .A(n37), .ZN(n253) );
  INV_X1 U273 ( .A(n41), .ZN(n260) );
  INV_X1 U274 ( .A(n185), .ZN(n266) );
  AOI22_X1 U275 ( .A1(b[54]), .A2(a[54]), .B1(n166), .B2(n81), .ZN(n138) );
  AOI22_X1 U276 ( .A1(b[34]), .A2(a[34]), .B1(n225), .B2(n103), .ZN(n158) );
  AOI22_X1 U277 ( .A1(b[24]), .A2(a[24]), .B1(n221), .B2(n114), .ZN(n168) );
  AOI22_X1 U278 ( .A1(b[14]), .A2(a[14]), .B1(n217), .B2(n125), .ZN(n178) );
  AOI22_X1 U279 ( .A1(b[60]), .A2(a[60]), .B1(n39), .B2(n74), .ZN(n132) );
  AOI22_X1 U280 ( .A1(b[32]), .A2(a[32]), .B1(n27), .B2(n105), .ZN(n160) );
  AOI22_X1 U281 ( .A1(b[22]), .A2(a[22]), .B1(n254), .B2(n116), .ZN(n170) );
  AOI22_X1 U282 ( .A1(b[12]), .A2(a[12]), .B1(n261), .B2(n127), .ZN(n180) );
  AOI22_X1 U283 ( .A1(b[5]), .A2(a[5]), .B1(n268), .B2(n75), .ZN(n186) );
  INV_X1 U284 ( .A(n187), .ZN(n268) );
  AOI22_X1 U285 ( .A1(b[6]), .A2(a[6]), .B1(n267), .B2(n69), .ZN(n185) );
  INV_X1 U286 ( .A(n186), .ZN(n267) );
  INV_X1 U287 ( .A(n1), .ZN(n232) );
  INV_X1 U288 ( .A(n35), .ZN(n235) );
  INV_X1 U289 ( .A(n2), .ZN(n244) );
  INV_X1 U290 ( .A(n131), .ZN(n249) );
  INV_X1 U291 ( .A(n40), .ZN(n256) );
  INV_X1 U292 ( .A(n191), .ZN(n272) );
  OAI22_X1 U293 ( .A1(n230), .A2(n273), .B1(n216), .B2(n70), .ZN(cout) );
  XNOR2_X1 U294 ( .A(n65), .B(n10), .ZN(result[9]) );
  INV_X1 U295 ( .A(n4), .ZN(n233) );
  INV_X1 U296 ( .A(n141), .ZN(n236) );
  INV_X1 U297 ( .A(n195), .ZN(n238) );
  INV_X1 U298 ( .A(n146), .ZN(n239) );
  INV_X1 U299 ( .A(n149), .ZN(n241) );
  INV_X1 U300 ( .A(n36), .ZN(n242) );
  INV_X1 U301 ( .A(n156), .ZN(n245) );
  INV_X1 U302 ( .A(n165), .ZN(n250) );
  INV_X1 U303 ( .A(n171), .ZN(n254) );
  INV_X1 U304 ( .A(n175), .ZN(n257) );
  INV_X1 U305 ( .A(n181), .ZN(n261) );
  AOI22_X1 U306 ( .A1(b[0]), .A2(a[0]), .B1(n130), .B2(cin), .ZN(n191) );
  INV_X1 U307 ( .A(n3), .ZN(n234) );
  AOI22_X1 U308 ( .A1(b[56]), .A2(a[56]), .B1(n53), .B2(n79), .ZN(n136) );
  INV_X1 U309 ( .A(n5), .ZN(n237) );
  AOI22_X1 U310 ( .A1(b[51]), .A2(a[51]), .B1(n31), .B2(n84), .ZN(n141) );
  AOI22_X1 U311 ( .A1(b[45]), .A2(a[45]), .B1(n23), .B2(n91), .ZN(n147) );
  AOI22_X1 U312 ( .A1(b[46]), .A2(a[46]), .B1(n240), .B2(n90), .ZN(n146) );
  INV_X1 U313 ( .A(n147), .ZN(n240) );
  AOI22_X1 U314 ( .A1(b[40]), .A2(a[40]), .B1(n57), .B2(n96), .ZN(n152) );
  AOI22_X1 U315 ( .A1(b[41]), .A2(a[41]), .B1(n243), .B2(n95), .ZN(n151) );
  INV_X1 U316 ( .A(n152), .ZN(n243) );
  INV_X1 U317 ( .A(n158), .ZN(n246) );
  AOI22_X1 U318 ( .A1(b[36]), .A2(a[36]), .B1(n49), .B2(n101), .ZN(n156) );
  AOI22_X1 U319 ( .A1(b[30]), .A2(a[30]), .B1(n137), .B2(n107), .ZN(n162) );
  INV_X1 U320 ( .A(n162), .ZN(n248) );
  AOI22_X1 U321 ( .A1(b[25]), .A2(a[25]), .B1(n252), .B2(n113), .ZN(n167) );
  INV_X1 U322 ( .A(n168), .ZN(n252) );
  INV_X1 U323 ( .A(n38), .ZN(n251) );
  AOI22_X1 U324 ( .A1(b[20]), .A2(a[20]), .B1(n208), .B2(n118), .ZN(n172) );
  AOI22_X1 U325 ( .A1(b[21]), .A2(a[21]), .B1(n255), .B2(n117), .ZN(n171) );
  INV_X1 U326 ( .A(n172), .ZN(n255) );
  AOI22_X1 U327 ( .A1(b[15]), .A2(a[15]), .B1(n259), .B2(n124), .ZN(n177) );
  INV_X1 U328 ( .A(n178), .ZN(n259) );
  INV_X1 U329 ( .A(n133), .ZN(n258) );
  AOI22_X1 U330 ( .A1(b[10]), .A2(a[10]), .B1(n263), .B2(n129), .ZN(n182) );
  INV_X1 U331 ( .A(n183), .ZN(n263) );
  AOI22_X1 U332 ( .A1(b[11]), .A2(a[11]), .B1(n262), .B2(n128), .ZN(n181) );
  INV_X1 U333 ( .A(n182), .ZN(n262) );
  AOI22_X1 U334 ( .A1(b[9]), .A2(a[9]), .B1(n264), .B2(n65), .ZN(n183) );
  INV_X1 U335 ( .A(n66), .ZN(n264) );
  AOI22_X1 U336 ( .A1(b[62]), .A2(a[62]), .B1(n45), .B2(n72), .ZN(n71) );
  AOI22_X1 U337 ( .A1(b[8]), .A2(a[8]), .B1(n265), .B2(n67), .ZN(n66) );
  INV_X1 U338 ( .A(n184), .ZN(n265) );
endmodule


module sequentialMultiplier ( a, b, reset, clk, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;
  input reset, clk;
  wire   N1, N2, N3, N4, N5, n_0_net__63_, n_0_net__62_, n_0_net__61_,
         n_0_net__60_, n_0_net__59_, n_0_net__58_, n_0_net__57_, n_0_net__56_,
         n_0_net__55_, n_0_net__54_, n_0_net__53_, n_0_net__52_, n_0_net__51_,
         n_0_net__50_, n_0_net__49_, n_0_net__48_, n_0_net__47_, n_0_net__46_,
         n_0_net__45_, n_0_net__44_, n_0_net__43_, n_0_net__42_, n_0_net__41_,
         n_0_net__40_, n_0_net__39_, n_0_net__38_, n_0_net__37_, n_0_net__36_,
         n_0_net__35_, n_0_net__34_, n_0_net__33_, n_0_net__32_, n_0_net__31_,
         n_0_net__30_, n_0_net__29_, n_0_net__28_, n_0_net__27_, n_0_net__26_,
         n_0_net__25_, n_0_net__24_, n_0_net__23_, n_0_net__22_, n_0_net__21_,
         n_0_net__20_, n_0_net__19_, n_0_net__18_, n_0_net__17_, n_0_net__16_,
         n_0_net__15_, n_0_net__14_, n_0_net__13_, n_0_net__12_, n_0_net__11_,
         n_0_net__10_, n_0_net__9_, n_0_net__8_, n_0_net__7_, n_0_net__6_,
         n_0_net__5_, n_0_net__4_, n_0_net__3_, n_0_net__2_, n_0_net__1_,
         n_0_net__0_, i_5_, N6, N7, N8, N9, N11, N12, N13, N14, N15, N16, N17,
         N18, N20, N21, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39,
         N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67,
         N68, N69, N74, N76, N77, N78, N79, N80, N146, N147, N148, N149, N150,
         N151, n67, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137,
         sll_14_ML_int_5__16_, sll_14_ML_int_5__17_, sll_14_ML_int_5__18_,
         sll_14_ML_int_5__19_, sll_14_ML_int_5__20_, sll_14_ML_int_5__21_,
         sll_14_ML_int_5__22_, sll_14_ML_int_5__23_, sll_14_ML_int_5__24_,
         sll_14_ML_int_5__25_, sll_14_ML_int_5__26_, sll_14_ML_int_5__27_,
         sll_14_ML_int_5__28_, sll_14_ML_int_5__29_, sll_14_ML_int_5__30_,
         sll_14_ML_int_5__31_, sll_14_ML_int_5__32_, sll_14_ML_int_5__33_,
         sll_14_ML_int_5__34_, sll_14_ML_int_5__35_, sll_14_ML_int_5__36_,
         sll_14_ML_int_5__37_, sll_14_ML_int_5__38_, sll_14_ML_int_5__39_,
         sll_14_ML_int_5__40_, sll_14_ML_int_5__41_, sll_14_ML_int_5__42_,
         sll_14_ML_int_5__43_, sll_14_ML_int_5__44_, sll_14_ML_int_5__45_,
         sll_14_ML_int_5__46_, sll_14_ML_int_5__47_, sll_14_ML_int_5__48_,
         sll_14_ML_int_5__49_, sll_14_ML_int_5__50_, sll_14_ML_int_5__51_,
         sll_14_ML_int_5__52_, sll_14_ML_int_5__53_, sll_14_ML_int_5__54_,
         sll_14_ML_int_5__55_, sll_14_ML_int_5__56_, sll_14_ML_int_5__57_,
         sll_14_ML_int_5__58_, sll_14_ML_int_5__59_, sll_14_ML_int_5__60_,
         sll_14_ML_int_5__61_, sll_14_ML_int_4__0_, sll_14_ML_int_4__1_,
         sll_14_ML_int_4__2_, sll_14_ML_int_4__3_, sll_14_ML_int_4__4_,
         sll_14_ML_int_4__5_, sll_14_ML_int_4__6_, sll_14_ML_int_4__7_,
         sll_14_ML_int_4__8_, sll_14_ML_int_4__9_, sll_14_ML_int_4__10_,
         sll_14_ML_int_4__11_, sll_14_ML_int_4__12_, sll_14_ML_int_4__13_,
         sll_14_ML_int_4__14_, sll_14_ML_int_4__15_, sll_14_ML_int_4__16_,
         sll_14_ML_int_4__17_, sll_14_ML_int_4__18_, sll_14_ML_int_4__19_,
         sll_14_ML_int_4__20_, sll_14_ML_int_4__21_, sll_14_ML_int_4__22_,
         sll_14_ML_int_4__23_, sll_14_ML_int_4__24_, sll_14_ML_int_4__25_,
         sll_14_ML_int_4__26_, sll_14_ML_int_4__27_, sll_14_ML_int_4__28_,
         sll_14_ML_int_4__29_, sll_14_ML_int_4__30_, sll_14_ML_int_4__32_,
         sll_14_ML_int_4__33_, sll_14_ML_int_4__34_, sll_14_ML_int_4__35_,
         sll_14_ML_int_4__36_, sll_14_ML_int_4__37_, sll_14_ML_int_4__38_,
         sll_14_ML_int_4__39_, sll_14_ML_int_4__40_, sll_14_ML_int_4__41_,
         sll_14_ML_int_4__42_, sll_14_ML_int_4__43_, sll_14_ML_int_4__44_,
         sll_14_ML_int_4__45_, sll_14_ML_int_3__1_, sll_14_ML_int_3__2_,
         sll_14_ML_int_3__3_, sll_14_ML_int_3__4_, sll_14_ML_int_3__5_,
         sll_14_ML_int_3__6_, sll_14_ML_int_3__7_, sll_14_ML_int_3__8_,
         sll_14_ML_int_3__9_, sll_14_ML_int_3__10_, sll_14_ML_int_3__11_,
         sll_14_ML_int_3__12_, sll_14_ML_int_3__13_, sll_14_ML_int_3__14_,
         sll_14_ML_int_3__15_, sll_14_ML_int_3__16_, sll_14_ML_int_3__17_,
         sll_14_ML_int_3__18_, sll_14_ML_int_3__19_, sll_14_ML_int_3__20_,
         sll_14_ML_int_3__21_, sll_14_ML_int_3__22_, sll_14_ML_int_3__23_,
         sll_14_ML_int_3__24_, sll_14_ML_int_3__25_, sll_14_ML_int_3__26_,
         sll_14_ML_int_3__27_, sll_14_ML_int_3__28_, sll_14_ML_int_3__29_,
         sll_14_ML_int_3__30_, sll_14_ML_int_2__0_, sll_14_ML_int_2__1_,
         sll_14_ML_int_2__2_, sll_14_ML_int_2__3_, sll_14_ML_int_2__4_,
         sll_14_ML_int_2__5_, sll_14_ML_int_2__6_, sll_14_ML_int_2__7_,
         sll_14_ML_int_2__8_, sll_14_ML_int_2__9_, sll_14_ML_int_2__10_,
         sll_14_ML_int_2__11_, sll_14_ML_int_2__12_, sll_14_ML_int_2__13_,
         sll_14_ML_int_2__14_, sll_14_ML_int_2__15_, sll_14_ML_int_2__16_,
         sll_14_ML_int_2__17_, sll_14_ML_int_2__18_, sll_14_ML_int_2__19_,
         sll_14_ML_int_2__20_, sll_14_ML_int_2__21_, sll_14_ML_int_2__22_,
         sll_14_ML_int_2__23_, sll_14_ML_int_2__24_, sll_14_ML_int_2__25_,
         sll_14_ML_int_2__26_, sll_14_ML_int_2__27_, sll_14_ML_int_2__28_,
         sll_14_ML_int_2__29_, sll_14_ML_int_2__30_, sll_14_ML_int_1__0_,
         sll_14_ML_int_1__1_, sll_14_ML_int_1__2_, sll_14_ML_int_1__3_,
         sll_14_ML_int_1__4_, sll_14_ML_int_1__5_, sll_14_ML_int_1__6_,
         sll_14_ML_int_1__7_, sll_14_ML_int_1__8_, sll_14_ML_int_1__9_,
         sll_14_ML_int_1__10_, sll_14_ML_int_1__11_, sll_14_ML_int_1__12_,
         sll_14_ML_int_1__13_, sll_14_ML_int_1__14_, sll_14_ML_int_1__15_,
         sll_14_ML_int_1__16_, sll_14_ML_int_1__17_, sll_14_ML_int_1__18_,
         sll_14_ML_int_1__19_, sll_14_ML_int_1__20_, sll_14_ML_int_1__21_,
         sll_14_ML_int_1__22_, sll_14_ML_int_1__23_, sll_14_ML_int_1__24_,
         sll_14_ML_int_1__25_, sll_14_ML_int_1__26_, sll_14_ML_int_1__27_,
         sll_14_ML_int_1__28_, sll_14_ML_int_1__29_, sll_14_ML_int_1__30_, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n68, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325;
  wire   [63:0] tempResult;
  wire   [5:2] add_30_carry;

  DFF_X1 i_reg_0_ ( .D(N146), .CK(clk), .Q(N1), .QN(n182) );
  DFF_X1 i_reg_5_ ( .D(N151), .CK(clk), .Q(i_5_), .QN(n67) );
  DFF_X1 i_reg_4_ ( .D(N150), .CK(clk), .Q(N5), .QN(n176) );
  DFF_X1 i_reg_3_ ( .D(N149), .CK(clk), .Q(N4), .QN(n177) );
  DFF_X1 i_reg_2_ ( .D(N148), .CK(clk), .Q(N3), .QN(n180) );
  DFF_X1 i_reg_1_ ( .D(N147), .CK(clk), .Q(N2), .QN(n181) );
  DFF_X1 A_reg_0_ ( .D(n324), .CK(clk), .Q(result[0]) );
  DFF_X1 A_reg_1_ ( .D(n323), .CK(clk), .Q(result[1]) );
  DFF_X1 A_reg_2_ ( .D(n322), .CK(clk), .Q(result[2]) );
  DFF_X1 A_reg_3_ ( .D(n321), .CK(clk), .Q(result[3]) );
  DFF_X1 A_reg_4_ ( .D(n320), .CK(clk), .Q(result[4]) );
  DFF_X1 A_reg_5_ ( .D(n319), .CK(clk), .Q(result[5]) );
  DFF_X1 A_reg_6_ ( .D(n318), .CK(clk), .Q(result[6]) );
  DFF_X1 A_reg_7_ ( .D(n317), .CK(clk), .Q(result[7]) );
  DFF_X1 A_reg_8_ ( .D(n316), .CK(clk), .Q(result[8]) );
  DFF_X1 A_reg_9_ ( .D(n315), .CK(clk), .Q(result[9]) );
  DFF_X1 A_reg_10_ ( .D(n314), .CK(clk), .Q(result[10]) );
  DFF_X1 A_reg_11_ ( .D(n313), .CK(clk), .Q(result[11]) );
  DFF_X1 A_reg_12_ ( .D(n312), .CK(clk), .Q(result[12]) );
  DFF_X1 A_reg_13_ ( .D(n311), .CK(clk), .Q(result[13]) );
  DFF_X1 A_reg_14_ ( .D(n310), .CK(clk), .Q(result[14]) );
  DFF_X1 A_reg_15_ ( .D(n309), .CK(clk), .Q(result[15]) );
  DFF_X1 A_reg_16_ ( .D(n308), .CK(clk), .Q(result[16]) );
  DFF_X1 A_reg_17_ ( .D(n307), .CK(clk), .Q(result[17]) );
  DFF_X1 A_reg_18_ ( .D(n306), .CK(clk), .Q(result[18]) );
  DFF_X1 A_reg_19_ ( .D(n305), .CK(clk), .Q(result[19]) );
  DFF_X1 A_reg_20_ ( .D(n304), .CK(clk), .Q(result[20]) );
  DFF_X1 A_reg_21_ ( .D(n303), .CK(clk), .Q(result[21]) );
  DFF_X1 A_reg_22_ ( .D(n302), .CK(clk), .Q(result[22]) );
  DFF_X1 A_reg_23_ ( .D(n301), .CK(clk), .Q(result[23]) );
  DFF_X1 A_reg_24_ ( .D(n300), .CK(clk), .Q(result[24]) );
  DFF_X1 A_reg_25_ ( .D(n299), .CK(clk), .Q(result[25]) );
  DFF_X1 A_reg_26_ ( .D(n298), .CK(clk), .Q(result[26]) );
  DFF_X1 A_reg_27_ ( .D(n297), .CK(clk), .Q(result[27]) );
  DFF_X1 A_reg_28_ ( .D(n296), .CK(clk), .Q(result[28]) );
  DFF_X1 A_reg_29_ ( .D(n295), .CK(clk), .Q(result[29]) );
  DFF_X1 A_reg_30_ ( .D(n294), .CK(clk), .Q(result[30]) );
  DFF_X1 A_reg_31_ ( .D(n293), .CK(clk), .Q(result[31]) );
  DFF_X1 A_reg_32_ ( .D(n292), .CK(clk), .Q(result[32]) );
  DFF_X1 A_reg_33_ ( .D(n291), .CK(clk), .Q(result[33]) );
  DFF_X1 A_reg_34_ ( .D(n290), .CK(clk), .Q(result[34]) );
  DFF_X1 A_reg_35_ ( .D(n289), .CK(clk), .Q(result[35]) );
  DFF_X1 A_reg_36_ ( .D(n288), .CK(clk), .Q(result[36]) );
  DFF_X1 A_reg_37_ ( .D(n287), .CK(clk), .Q(result[37]) );
  DFF_X1 A_reg_38_ ( .D(n286), .CK(clk), .Q(result[38]) );
  DFF_X1 A_reg_39_ ( .D(n285), .CK(clk), .Q(result[39]) );
  DFF_X1 A_reg_40_ ( .D(n284), .CK(clk), .Q(result[40]) );
  DFF_X1 A_reg_41_ ( .D(n283), .CK(clk), .Q(result[41]) );
  DFF_X1 A_reg_42_ ( .D(n282), .CK(clk), .Q(result[42]) );
  DFF_X1 A_reg_43_ ( .D(n281), .CK(clk), .Q(result[43]) );
  DFF_X1 A_reg_44_ ( .D(n280), .CK(clk), .Q(result[44]) );
  DFF_X1 A_reg_45_ ( .D(n279), .CK(clk), .Q(result[45]) );
  DFF_X1 A_reg_46_ ( .D(n278), .CK(clk), .Q(result[46]) );
  DFF_X1 A_reg_47_ ( .D(n277), .CK(clk), .Q(result[47]) );
  DFF_X1 A_reg_48_ ( .D(n276), .CK(clk), .Q(result[48]) );
  DFF_X1 A_reg_49_ ( .D(n275), .CK(clk), .Q(result[49]) );
  DFF_X1 A_reg_50_ ( .D(n274), .CK(clk), .Q(result[50]) );
  DFF_X1 A_reg_51_ ( .D(n273), .CK(clk), .Q(result[51]) );
  DFF_X1 A_reg_52_ ( .D(n272), .CK(clk), .Q(result[52]) );
  DFF_X1 A_reg_53_ ( .D(n271), .CK(clk), .Q(result[53]) );
  DFF_X1 A_reg_54_ ( .D(n270), .CK(clk), .Q(result[54]) );
  DFF_X1 A_reg_55_ ( .D(n269), .CK(clk), .Q(result[55]) );
  DFF_X1 A_reg_56_ ( .D(n268), .CK(clk), .Q(result[56]) );
  DFF_X1 A_reg_57_ ( .D(n267), .CK(clk), .Q(result[57]) );
  DFF_X1 A_reg_58_ ( .D(n266), .CK(clk), .Q(result[58]) );
  DFF_X1 A_reg_59_ ( .D(n265), .CK(clk), .Q(result[59]) );
  DFF_X1 A_reg_60_ ( .D(n264), .CK(clk), .Q(result[60]) );
  DFF_X1 A_reg_61_ ( .D(n263), .CK(clk), .Q(result[61]) );
  DFF_X1 A_reg_62_ ( .D(n262), .CK(clk), .Q(result[62]) );
  XOR2_X1 U144 ( .A(N15), .B(n152), .Z(n_0_net__9_) );
  XOR2_X1 U145 ( .A(N14), .B(n150), .Z(n_0_net__8_) );
  XOR2_X1 U146 ( .A(N13), .B(n149), .Z(n_0_net__7_) );
  XOR2_X1 U147 ( .A(N12), .B(n148), .Z(n_0_net__6_) );
  XOR2_X1 U148 ( .A(N69), .B(n174), .Z(n_0_net__63_) );
  XOR2_X1 U149 ( .A(N68), .B(n173), .Z(n_0_net__62_) );
  XOR2_X1 U150 ( .A(N67), .B(n172), .Z(n_0_net__61_) );
  XOR2_X1 U151 ( .A(N66), .B(n171), .Z(n_0_net__60_) );
  XOR2_X1 U152 ( .A(N11), .B(n147), .Z(n_0_net__5_) );
  XOR2_X1 U153 ( .A(N65), .B(n170), .Z(n_0_net__59_) );
  XOR2_X1 U154 ( .A(N64), .B(n167), .Z(n_0_net__58_) );
  XOR2_X1 U155 ( .A(N63), .B(n166), .Z(n_0_net__57_) );
  XOR2_X1 U156 ( .A(N62), .B(n165), .Z(n_0_net__56_) );
  XOR2_X1 U158 ( .A(N60), .B(n163), .Z(n_0_net__54_) );
  XOR2_X1 U159 ( .A(N59), .B(n162), .Z(n_0_net__53_) );
  XOR2_X1 U160 ( .A(N58), .B(n161), .Z(n_0_net__52_) );
  XOR2_X1 U161 ( .A(N57), .B(n160), .Z(n_0_net__51_) );
  XOR2_X1 U164 ( .A(N55), .B(n158), .Z(n_0_net__49_) );
  XOR2_X1 U166 ( .A(N53), .B(n156), .Z(n_0_net__47_) );
  XOR2_X1 U167 ( .A(N52), .B(n152), .Z(n_0_net__46_) );
  XOR2_X1 U168 ( .A(N51), .B(n151), .Z(n_0_net__45_) );
  XOR2_X1 U170 ( .A(N49), .B(n149), .Z(n_0_net__43_) );
  XOR2_X1 U172 ( .A(N47), .B(n147), .Z(n_0_net__41_) );
  XOR2_X1 U173 ( .A(N46), .B(n146), .Z(n_0_net__40_) );
  XOR2_X1 U174 ( .A(N9), .B(n145), .Z(n_0_net__3_) );
  XOR2_X1 U175 ( .A(N45), .B(n145), .Z(n_0_net__39_) );
  XOR2_X1 U176 ( .A(N44), .B(n144), .Z(n_0_net__38_) );
  XOR2_X1 U177 ( .A(N43), .B(n143), .Z(n_0_net__37_) );
  XOR2_X1 U178 ( .A(N42), .B(n142), .Z(n_0_net__36_) );
  XOR2_X1 U179 ( .A(N41), .B(n142), .Z(n_0_net__35_) );
  XOR2_X1 U181 ( .A(N39), .B(n171), .Z(n_0_net__33_) );
  XOR2_X1 U183 ( .A(N37), .B(n175), .Z(n_0_net__31_) );
  XOR2_X1 U184 ( .A(N36), .B(n175), .Z(n_0_net__30_) );
  XOR2_X1 U185 ( .A(N8), .B(n144), .Z(n_0_net__2_) );
  XOR2_X1 U186 ( .A(N35), .B(n142), .Z(n_0_net__29_) );
  XOR2_X1 U187 ( .A(N34), .B(n175), .Z(n_0_net__28_) );
  XOR2_X1 U188 ( .A(N33), .B(n171), .Z(n_0_net__27_) );
  XOR2_X1 U190 ( .A(N31), .B(n173), .Z(n_0_net__25_) );
  XOR2_X1 U191 ( .A(N30), .B(n172), .Z(n_0_net__24_) );
  XOR2_X1 U192 ( .A(N29), .B(n159), .Z(n_0_net__23_) );
  XOR2_X1 U196 ( .A(N7), .B(n137), .Z(n_0_net__1_) );
  XOR2_X1 U201 ( .A(N21), .B(n161), .Z(n_0_net__15_) );
  XOR2_X1 U202 ( .A(N20), .B(n160), .Z(n_0_net__14_) );
  XOR2_X1 U204 ( .A(N18), .B(n158), .Z(n_0_net__12_) );
  XOR2_X1 U205 ( .A(N17), .B(n157), .Z(n_0_net__11_) );
  XOR2_X1 U206 ( .A(N16), .B(n156), .Z(n_0_net__10_) );
  carryLookAheadAdder64bit A0 ( .a(result), .b({n_0_net__63_, n_0_net__62_, 
        n_0_net__61_, n_0_net__60_, n_0_net__59_, n_0_net__58_, n_0_net__57_, 
        n_0_net__56_, n_0_net__55_, n_0_net__54_, n_0_net__53_, n_0_net__52_, 
        n_0_net__51_, n_0_net__50_, n_0_net__49_, n_0_net__48_, n_0_net__47_, 
        n_0_net__46_, n_0_net__45_, n_0_net__44_, n_0_net__43_, n_0_net__42_, 
        n_0_net__41_, n_0_net__40_, n_0_net__39_, n_0_net__38_, n_0_net__37_, 
        n_0_net__36_, n_0_net__35_, n_0_net__34_, n_0_net__33_, n_0_net__32_, 
        n_0_net__31_, n_0_net__30_, n_0_net__29_, n_0_net__28_, n_0_net__27_, 
        n_0_net__26_, n_0_net__25_, n_0_net__24_, n_0_net__23_, n_0_net__22_, 
        n_0_net__21_, n_0_net__20_, n_0_net__19_, n_0_net__18_, n_0_net__17_, 
        n_0_net__16_, n_0_net__15_, n_0_net__14_, n_0_net__13_, n_0_net__12_, 
        n_0_net__11_, n_0_net__10_, n_0_net__9_, n_0_net__8_, n_0_net__7_, 
        n_0_net__6_, n_0_net__5_, n_0_net__4_, n_0_net__3_, n_0_net__2_, 
        n_0_net__1_, n_0_net__0_}), .cin(n143), .result(tempResult) );
  HA_X1 add_30_U1_1_1 ( .A(n215), .B(n66), .CO(add_30_carry[2]), .S(N76) );
  HA_X1 add_30_U1_1_2 ( .A(n213), .B(add_30_carry[2]), .CO(add_30_carry[3]), 
        .S(N77) );
  HA_X1 add_30_U1_1_3 ( .A(n209), .B(add_30_carry[3]), .CO(add_30_carry[4]), 
        .S(N78) );
  HA_X1 add_30_U1_1_4 ( .A(n206), .B(add_30_carry[4]), .CO(add_30_carry[5]), 
        .S(N79) );
  MUX2_X1 sll_14_M1_0_1 ( .A(a[1]), .B(a[0]), .S(N1), .Z(sll_14_ML_int_1__1_)
         );
  MUX2_X1 sll_14_M1_0_3 ( .A(a[3]), .B(a[2]), .S(n217), .Z(sll_14_ML_int_1__3_) );
  MUX2_X1 sll_14_M1_0_4 ( .A(a[4]), .B(a[3]), .S(n217), .Z(sll_14_ML_int_1__4_) );
  MUX2_X1 sll_14_M1_0_5 ( .A(a[5]), .B(a[4]), .S(n12), .Z(sll_14_ML_int_1__5_)
         );
  MUX2_X1 sll_14_M1_0_6 ( .A(a[6]), .B(a[5]), .S(n12), .Z(sll_14_ML_int_1__6_)
         );
  MUX2_X1 sll_14_M1_0_7 ( .A(a[7]), .B(a[6]), .S(n12), .Z(sll_14_ML_int_1__7_)
         );
  MUX2_X1 sll_14_M1_0_8 ( .A(a[8]), .B(a[7]), .S(n12), .Z(sll_14_ML_int_1__8_)
         );
  MUX2_X1 sll_14_M1_0_9 ( .A(a[9]), .B(a[8]), .S(n12), .Z(sll_14_ML_int_1__9_)
         );
  MUX2_X1 sll_14_M1_0_10 ( .A(a[10]), .B(a[9]), .S(n12), .Z(
        sll_14_ML_int_1__10_) );
  MUX2_X1 sll_14_M1_0_11 ( .A(a[11]), .B(a[10]), .S(n12), .Z(
        sll_14_ML_int_1__11_) );
  MUX2_X1 sll_14_M1_0_12 ( .A(a[12]), .B(a[11]), .S(n12), .Z(
        sll_14_ML_int_1__12_) );
  MUX2_X1 sll_14_M1_0_13 ( .A(a[13]), .B(a[12]), .S(n12), .Z(
        sll_14_ML_int_1__13_) );
  MUX2_X1 sll_14_M1_0_14 ( .A(a[14]), .B(a[13]), .S(n12), .Z(
        sll_14_ML_int_1__14_) );
  MUX2_X1 sll_14_M1_0_15 ( .A(a[15]), .B(a[14]), .S(n12), .Z(
        sll_14_ML_int_1__15_) );
  MUX2_X1 sll_14_M1_0_16 ( .A(a[16]), .B(a[15]), .S(n12), .Z(
        sll_14_ML_int_1__16_) );
  MUX2_X1 sll_14_M1_0_17 ( .A(a[17]), .B(a[16]), .S(n12), .Z(
        sll_14_ML_int_1__17_) );
  MUX2_X1 sll_14_M1_0_18 ( .A(a[18]), .B(a[17]), .S(n66), .Z(
        sll_14_ML_int_1__18_) );
  MUX2_X1 sll_14_M1_0_19 ( .A(a[19]), .B(a[18]), .S(n12), .Z(
        sll_14_ML_int_1__19_) );
  MUX2_X1 sll_14_M1_0_20 ( .A(a[20]), .B(a[19]), .S(n66), .Z(
        sll_14_ML_int_1__20_) );
  MUX2_X1 sll_14_M1_0_21 ( .A(a[21]), .B(a[20]), .S(n66), .Z(
        sll_14_ML_int_1__21_) );
  MUX2_X1 sll_14_M1_0_22 ( .A(a[22]), .B(a[21]), .S(n66), .Z(
        sll_14_ML_int_1__22_) );
  MUX2_X1 sll_14_M1_0_23 ( .A(a[23]), .B(a[22]), .S(n66), .Z(
        sll_14_ML_int_1__23_) );
  MUX2_X1 sll_14_M1_0_24 ( .A(a[24]), .B(a[23]), .S(n66), .Z(
        sll_14_ML_int_1__24_) );
  MUX2_X1 sll_14_M1_0_25 ( .A(a[25]), .B(a[24]), .S(n66), .Z(
        sll_14_ML_int_1__25_) );
  MUX2_X1 sll_14_M1_0_26 ( .A(a[26]), .B(a[25]), .S(n66), .Z(
        sll_14_ML_int_1__26_) );
  MUX2_X1 sll_14_M1_0_27 ( .A(a[27]), .B(a[26]), .S(n66), .Z(
        sll_14_ML_int_1__27_) );
  MUX2_X1 sll_14_M1_0_28 ( .A(a[28]), .B(a[27]), .S(n66), .Z(
        sll_14_ML_int_1__28_) );
  MUX2_X1 sll_14_M1_0_29 ( .A(a[29]), .B(a[28]), .S(n66), .Z(
        sll_14_ML_int_1__29_) );
  MUX2_X1 sll_14_M1_0_30 ( .A(a[30]), .B(a[29]), .S(n66), .Z(
        sll_14_ML_int_1__30_) );
  MUX2_X1 sll_14_M1_1_4 ( .A(sll_14_ML_int_1__4_), .B(n11), .S(n216), .Z(
        sll_14_ML_int_2__4_) );
  MUX2_X1 sll_14_M1_1_5 ( .A(sll_14_ML_int_1__5_), .B(sll_14_ML_int_1__3_), 
        .S(n215), .Z(sll_14_ML_int_2__5_) );
  MUX2_X1 sll_14_M1_1_6 ( .A(sll_14_ML_int_1__6_), .B(sll_14_ML_int_1__4_), 
        .S(n215), .Z(sll_14_ML_int_2__6_) );
  MUX2_X1 sll_14_M1_1_7 ( .A(sll_14_ML_int_1__7_), .B(sll_14_ML_int_1__5_), 
        .S(n215), .Z(sll_14_ML_int_2__7_) );
  MUX2_X1 sll_14_M1_1_8 ( .A(sll_14_ML_int_1__8_), .B(sll_14_ML_int_1__6_), 
        .S(n215), .Z(sll_14_ML_int_2__8_) );
  MUX2_X1 sll_14_M1_1_9 ( .A(sll_14_ML_int_1__9_), .B(sll_14_ML_int_1__7_), 
        .S(n215), .Z(sll_14_ML_int_2__9_) );
  MUX2_X1 sll_14_M1_1_10 ( .A(sll_14_ML_int_1__10_), .B(sll_14_ML_int_1__8_), 
        .S(n215), .Z(sll_14_ML_int_2__10_) );
  MUX2_X1 sll_14_M1_1_11 ( .A(sll_14_ML_int_1__11_), .B(sll_14_ML_int_1__9_), 
        .S(n215), .Z(sll_14_ML_int_2__11_) );
  MUX2_X1 sll_14_M1_1_12 ( .A(sll_14_ML_int_1__12_), .B(sll_14_ML_int_1__10_), 
        .S(n215), .Z(sll_14_ML_int_2__12_) );
  MUX2_X1 sll_14_M1_1_13 ( .A(sll_14_ML_int_1__13_), .B(sll_14_ML_int_1__11_), 
        .S(n215), .Z(sll_14_ML_int_2__13_) );
  MUX2_X1 sll_14_M1_1_14 ( .A(sll_14_ML_int_1__14_), .B(sll_14_ML_int_1__12_), 
        .S(n215), .Z(sll_14_ML_int_2__14_) );
  MUX2_X1 sll_14_M1_1_15 ( .A(sll_14_ML_int_1__15_), .B(sll_14_ML_int_1__13_), 
        .S(n215), .Z(sll_14_ML_int_2__15_) );
  MUX2_X1 sll_14_M1_1_16 ( .A(sll_14_ML_int_1__16_), .B(sll_14_ML_int_1__14_), 
        .S(n215), .Z(sll_14_ML_int_2__16_) );
  MUX2_X1 sll_14_M1_1_17 ( .A(sll_14_ML_int_1__17_), .B(sll_14_ML_int_1__15_), 
        .S(n215), .Z(sll_14_ML_int_2__17_) );
  MUX2_X1 sll_14_M1_1_18 ( .A(sll_14_ML_int_1__18_), .B(sll_14_ML_int_1__16_), 
        .S(n215), .Z(sll_14_ML_int_2__18_) );
  MUX2_X1 sll_14_M1_1_19 ( .A(sll_14_ML_int_1__19_), .B(sll_14_ML_int_1__17_), 
        .S(n215), .Z(sll_14_ML_int_2__19_) );
  MUX2_X1 sll_14_M1_1_20 ( .A(sll_14_ML_int_1__20_), .B(sll_14_ML_int_1__18_), 
        .S(n215), .Z(sll_14_ML_int_2__20_) );
  MUX2_X1 sll_14_M1_1_21 ( .A(sll_14_ML_int_1__21_), .B(sll_14_ML_int_1__19_), 
        .S(n215), .Z(sll_14_ML_int_2__21_) );
  MUX2_X1 sll_14_M1_1_22 ( .A(sll_14_ML_int_1__22_), .B(sll_14_ML_int_1__20_), 
        .S(n215), .Z(sll_14_ML_int_2__22_) );
  MUX2_X1 sll_14_M1_1_23 ( .A(sll_14_ML_int_1__23_), .B(sll_14_ML_int_1__21_), 
        .S(n215), .Z(sll_14_ML_int_2__23_) );
  MUX2_X1 sll_14_M1_1_24 ( .A(sll_14_ML_int_1__24_), .B(sll_14_ML_int_1__22_), 
        .S(n215), .Z(sll_14_ML_int_2__24_) );
  MUX2_X1 sll_14_M1_1_25 ( .A(sll_14_ML_int_1__25_), .B(sll_14_ML_int_1__23_), 
        .S(n215), .Z(sll_14_ML_int_2__25_) );
  MUX2_X1 sll_14_M1_1_26 ( .A(sll_14_ML_int_1__26_), .B(sll_14_ML_int_1__24_), 
        .S(n215), .Z(sll_14_ML_int_2__26_) );
  MUX2_X1 sll_14_M1_1_27 ( .A(sll_14_ML_int_1__27_), .B(sll_14_ML_int_1__25_), 
        .S(n216), .Z(sll_14_ML_int_2__27_) );
  MUX2_X1 sll_14_M1_1_28 ( .A(sll_14_ML_int_1__28_), .B(sll_14_ML_int_1__26_), 
        .S(n215), .Z(sll_14_ML_int_2__28_) );
  MUX2_X1 sll_14_M1_1_29 ( .A(sll_14_ML_int_1__29_), .B(sll_14_ML_int_1__27_), 
        .S(n215), .Z(sll_14_ML_int_2__29_) );
  MUX2_X1 sll_14_M1_1_30 ( .A(sll_14_ML_int_1__30_), .B(sll_14_ML_int_1__28_), 
        .S(n215), .Z(sll_14_ML_int_2__30_) );
  MUX2_X1 sll_14_M1_2_5 ( .A(sll_14_ML_int_2__5_), .B(n6), .S(n213), .Z(
        sll_14_ML_int_3__5_) );
  MUX2_X1 sll_14_M1_2_6 ( .A(sll_14_ML_int_2__6_), .B(n9), .S(n213), .Z(
        sll_14_ML_int_3__6_) );
  MUX2_X1 sll_14_M1_2_7 ( .A(sll_14_ML_int_2__7_), .B(sll_14_ML_int_2__3_), 
        .S(n213), .Z(sll_14_ML_int_3__7_) );
  MUX2_X1 sll_14_M1_2_8 ( .A(sll_14_ML_int_2__8_), .B(sll_14_ML_int_2__4_), 
        .S(n213), .Z(sll_14_ML_int_3__8_) );
  MUX2_X1 sll_14_M1_2_9 ( .A(sll_14_ML_int_2__9_), .B(sll_14_ML_int_2__5_), 
        .S(n213), .Z(sll_14_ML_int_3__9_) );
  MUX2_X1 sll_14_M1_2_10 ( .A(sll_14_ML_int_2__10_), .B(sll_14_ML_int_2__6_), 
        .S(n213), .Z(sll_14_ML_int_3__10_) );
  MUX2_X1 sll_14_M1_2_11 ( .A(sll_14_ML_int_2__11_), .B(sll_14_ML_int_2__7_), 
        .S(n213), .Z(sll_14_ML_int_3__11_) );
  MUX2_X1 sll_14_M1_2_12 ( .A(sll_14_ML_int_2__12_), .B(sll_14_ML_int_2__8_), 
        .S(n213), .Z(sll_14_ML_int_3__12_) );
  MUX2_X1 sll_14_M1_2_13 ( .A(sll_14_ML_int_2__13_), .B(sll_14_ML_int_2__9_), 
        .S(n213), .Z(sll_14_ML_int_3__13_) );
  MUX2_X1 sll_14_M1_2_14 ( .A(sll_14_ML_int_2__14_), .B(sll_14_ML_int_2__10_), 
        .S(n213), .Z(sll_14_ML_int_3__14_) );
  MUX2_X1 sll_14_M1_2_15 ( .A(sll_14_ML_int_2__15_), .B(sll_14_ML_int_2__11_), 
        .S(n213), .Z(sll_14_ML_int_3__15_) );
  MUX2_X1 sll_14_M1_2_16 ( .A(sll_14_ML_int_2__16_), .B(sll_14_ML_int_2__12_), 
        .S(n213), .Z(sll_14_ML_int_3__16_) );
  MUX2_X1 sll_14_M1_2_17 ( .A(sll_14_ML_int_2__17_), .B(sll_14_ML_int_2__13_), 
        .S(n213), .Z(sll_14_ML_int_3__17_) );
  MUX2_X1 sll_14_M1_2_18 ( .A(sll_14_ML_int_2__18_), .B(sll_14_ML_int_2__14_), 
        .S(n213), .Z(sll_14_ML_int_3__18_) );
  MUX2_X1 sll_14_M1_2_19 ( .A(sll_14_ML_int_2__19_), .B(sll_14_ML_int_2__15_), 
        .S(n213), .Z(sll_14_ML_int_3__19_) );
  MUX2_X1 sll_14_M1_2_20 ( .A(sll_14_ML_int_2__20_), .B(sll_14_ML_int_2__16_), 
        .S(n213), .Z(sll_14_ML_int_3__20_) );
  MUX2_X1 sll_14_M1_2_21 ( .A(sll_14_ML_int_2__21_), .B(sll_14_ML_int_2__17_), 
        .S(n213), .Z(sll_14_ML_int_3__21_) );
  MUX2_X1 sll_14_M1_2_22 ( .A(sll_14_ML_int_2__22_), .B(sll_14_ML_int_2__18_), 
        .S(n213), .Z(sll_14_ML_int_3__22_) );
  MUX2_X1 sll_14_M1_2_23 ( .A(sll_14_ML_int_2__23_), .B(sll_14_ML_int_2__19_), 
        .S(n213), .Z(sll_14_ML_int_3__23_) );
  MUX2_X1 sll_14_M1_2_24 ( .A(sll_14_ML_int_2__24_), .B(sll_14_ML_int_2__20_), 
        .S(n213), .Z(sll_14_ML_int_3__24_) );
  MUX2_X1 sll_14_M1_2_25 ( .A(sll_14_ML_int_2__25_), .B(sll_14_ML_int_2__21_), 
        .S(n213), .Z(sll_14_ML_int_3__25_) );
  MUX2_X1 sll_14_M1_2_26 ( .A(sll_14_ML_int_2__26_), .B(sll_14_ML_int_2__22_), 
        .S(n213), .Z(sll_14_ML_int_3__26_) );
  MUX2_X1 sll_14_M1_2_27 ( .A(sll_14_ML_int_2__27_), .B(sll_14_ML_int_2__23_), 
        .S(n213), .Z(sll_14_ML_int_3__27_) );
  MUX2_X1 sll_14_M1_2_28 ( .A(sll_14_ML_int_2__28_), .B(sll_14_ML_int_2__24_), 
        .S(n213), .Z(sll_14_ML_int_3__28_) );
  MUX2_X1 sll_14_M1_2_29 ( .A(sll_14_ML_int_2__29_), .B(sll_14_ML_int_2__25_), 
        .S(n213), .Z(sll_14_ML_int_3__29_) );
  MUX2_X1 sll_14_M1_2_30 ( .A(sll_14_ML_int_2__30_), .B(sll_14_ML_int_2__26_), 
        .S(n213), .Z(sll_14_ML_int_3__30_) );
  MUX2_X1 sll_14_M1_3_8 ( .A(sll_14_ML_int_3__8_), .B(n22), .S(n209), .Z(
        sll_14_ML_int_4__8_) );
  MUX2_X1 sll_14_M1_3_9 ( .A(sll_14_ML_int_3__9_), .B(sll_14_ML_int_3__1_), 
        .S(n209), .Z(sll_14_ML_int_4__9_) );
  MUX2_X1 sll_14_M1_3_10 ( .A(sll_14_ML_int_3__10_), .B(sll_14_ML_int_3__2_), 
        .S(n209), .Z(sll_14_ML_int_4__10_) );
  MUX2_X1 sll_14_M1_3_11 ( .A(sll_14_ML_int_3__11_), .B(sll_14_ML_int_3__3_), 
        .S(n209), .Z(sll_14_ML_int_4__11_) );
  MUX2_X1 sll_14_M1_3_12 ( .A(sll_14_ML_int_3__12_), .B(sll_14_ML_int_3__4_), 
        .S(n209), .Z(sll_14_ML_int_4__12_) );
  MUX2_X1 sll_14_M1_3_13 ( .A(sll_14_ML_int_3__13_), .B(sll_14_ML_int_3__5_), 
        .S(n209), .Z(sll_14_ML_int_4__13_) );
  MUX2_X1 sll_14_M1_3_14 ( .A(sll_14_ML_int_3__14_), .B(sll_14_ML_int_3__6_), 
        .S(n209), .Z(sll_14_ML_int_4__14_) );
  MUX2_X1 sll_14_M1_3_15 ( .A(sll_14_ML_int_3__15_), .B(sll_14_ML_int_3__7_), 
        .S(n209), .Z(sll_14_ML_int_4__15_) );
  MUX2_X1 sll_14_M1_3_16 ( .A(sll_14_ML_int_3__16_), .B(sll_14_ML_int_3__8_), 
        .S(n209), .Z(sll_14_ML_int_4__16_) );
  MUX2_X1 sll_14_M1_3_17 ( .A(sll_14_ML_int_3__17_), .B(sll_14_ML_int_3__9_), 
        .S(n209), .Z(sll_14_ML_int_4__17_) );
  MUX2_X1 sll_14_M1_3_18 ( .A(sll_14_ML_int_3__18_), .B(sll_14_ML_int_3__10_), 
        .S(n209), .Z(sll_14_ML_int_4__18_) );
  MUX2_X1 sll_14_M1_3_19 ( .A(sll_14_ML_int_3__19_), .B(sll_14_ML_int_3__11_), 
        .S(n210), .Z(sll_14_ML_int_4__19_) );
  MUX2_X1 sll_14_M1_3_20 ( .A(sll_14_ML_int_3__20_), .B(sll_14_ML_int_3__12_), 
        .S(n210), .Z(sll_14_ML_int_4__20_) );
  MUX2_X1 sll_14_M1_3_21 ( .A(sll_14_ML_int_3__21_), .B(sll_14_ML_int_3__13_), 
        .S(n210), .Z(sll_14_ML_int_4__21_) );
  MUX2_X1 sll_14_M1_3_22 ( .A(sll_14_ML_int_3__22_), .B(sll_14_ML_int_3__14_), 
        .S(n210), .Z(sll_14_ML_int_4__22_) );
  MUX2_X1 sll_14_M1_3_23 ( .A(sll_14_ML_int_3__23_), .B(sll_14_ML_int_3__15_), 
        .S(n210), .Z(sll_14_ML_int_4__23_) );
  MUX2_X1 sll_14_M1_3_24 ( .A(sll_14_ML_int_3__24_), .B(sll_14_ML_int_3__16_), 
        .S(n210), .Z(sll_14_ML_int_4__24_) );
  MUX2_X1 sll_14_M1_3_25 ( .A(sll_14_ML_int_3__25_), .B(sll_14_ML_int_3__17_), 
        .S(n210), .Z(sll_14_ML_int_4__25_) );
  MUX2_X1 sll_14_M1_3_26 ( .A(sll_14_ML_int_3__26_), .B(sll_14_ML_int_3__18_), 
        .S(n210), .Z(sll_14_ML_int_4__26_) );
  MUX2_X1 sll_14_M1_3_27 ( .A(sll_14_ML_int_3__27_), .B(sll_14_ML_int_3__19_), 
        .S(n210), .Z(sll_14_ML_int_4__27_) );
  MUX2_X1 sll_14_M1_3_28 ( .A(sll_14_ML_int_3__28_), .B(sll_14_ML_int_3__20_), 
        .S(n210), .Z(sll_14_ML_int_4__28_) );
  MUX2_X1 sll_14_M1_3_29 ( .A(sll_14_ML_int_3__29_), .B(sll_14_ML_int_3__21_), 
        .S(n210), .Z(sll_14_ML_int_4__29_) );
  MUX2_X1 sll_14_M1_3_30 ( .A(sll_14_ML_int_3__30_), .B(sll_14_ML_int_3__22_), 
        .S(n210), .Z(sll_14_ML_int_4__30_) );
  MUX2_X1 sll_14_M1_4_16 ( .A(sll_14_ML_int_4__16_), .B(sll_14_ML_int_4__0_), 
        .S(n206), .Z(sll_14_ML_int_5__16_) );
  MUX2_X1 sll_14_M1_4_17 ( .A(sll_14_ML_int_4__17_), .B(sll_14_ML_int_4__1_), 
        .S(n204), .Z(sll_14_ML_int_5__17_) );
  MUX2_X1 sll_14_M1_4_18 ( .A(sll_14_ML_int_4__18_), .B(sll_14_ML_int_4__2_), 
        .S(n204), .Z(sll_14_ML_int_5__18_) );
  MUX2_X1 sll_14_M1_4_19 ( .A(sll_14_ML_int_4__19_), .B(sll_14_ML_int_4__3_), 
        .S(n205), .Z(sll_14_ML_int_5__19_) );
  MUX2_X1 sll_14_M1_4_20 ( .A(sll_14_ML_int_4__20_), .B(sll_14_ML_int_4__4_), 
        .S(n204), .Z(sll_14_ML_int_5__20_) );
  MUX2_X1 sll_14_M1_4_21 ( .A(sll_14_ML_int_4__21_), .B(sll_14_ML_int_4__5_), 
        .S(n204), .Z(sll_14_ML_int_5__21_) );
  MUX2_X1 sll_14_M1_4_22 ( .A(sll_14_ML_int_4__22_), .B(sll_14_ML_int_4__6_), 
        .S(n204), .Z(sll_14_ML_int_5__22_) );
  MUX2_X1 sll_14_M1_4_23 ( .A(sll_14_ML_int_4__23_), .B(sll_14_ML_int_4__7_), 
        .S(n204), .Z(sll_14_ML_int_5__23_) );
  MUX2_X1 sll_14_M1_4_24 ( .A(sll_14_ML_int_4__24_), .B(sll_14_ML_int_4__8_), 
        .S(n204), .Z(sll_14_ML_int_5__24_) );
  MUX2_X1 sll_14_M1_4_25 ( .A(sll_14_ML_int_4__25_), .B(sll_14_ML_int_4__9_), 
        .S(n204), .Z(sll_14_ML_int_5__25_) );
  MUX2_X1 sll_14_M1_4_26 ( .A(sll_14_ML_int_4__26_), .B(sll_14_ML_int_4__10_), 
        .S(n204), .Z(sll_14_ML_int_5__26_) );
  MUX2_X1 sll_14_M1_4_27 ( .A(sll_14_ML_int_4__27_), .B(sll_14_ML_int_4__11_), 
        .S(n204), .Z(sll_14_ML_int_5__27_) );
  MUX2_X1 sll_14_M1_4_28 ( .A(sll_14_ML_int_4__28_), .B(sll_14_ML_int_4__12_), 
        .S(n204), .Z(sll_14_ML_int_5__28_) );
  MUX2_X1 sll_14_M1_4_29 ( .A(sll_14_ML_int_4__29_), .B(sll_14_ML_int_4__13_), 
        .S(n204), .Z(sll_14_ML_int_5__29_) );
  MUX2_X1 sll_14_M1_4_30 ( .A(sll_14_ML_int_4__30_), .B(sll_14_ML_int_4__14_), 
        .S(n204), .Z(sll_14_ML_int_5__30_) );
  MUX2_X1 sll_14_M1_4_32 ( .A(sll_14_ML_int_4__32_), .B(sll_14_ML_int_4__16_), 
        .S(n204), .Z(sll_14_ML_int_5__32_) );
  MUX2_X1 sll_14_M1_4_33 ( .A(sll_14_ML_int_4__33_), .B(sll_14_ML_int_4__17_), 
        .S(n206), .Z(sll_14_ML_int_5__33_) );
  MUX2_X1 sll_14_M1_4_34 ( .A(sll_14_ML_int_4__34_), .B(sll_14_ML_int_4__18_), 
        .S(n204), .Z(sll_14_ML_int_5__34_) );
  MUX2_X1 sll_14_M1_4_35 ( .A(sll_14_ML_int_4__35_), .B(sll_14_ML_int_4__19_), 
        .S(n204), .Z(sll_14_ML_int_5__35_) );
  MUX2_X1 sll_14_M1_4_36 ( .A(sll_14_ML_int_4__36_), .B(sll_14_ML_int_4__20_), 
        .S(n204), .Z(sll_14_ML_int_5__36_) );
  MUX2_X1 sll_14_M1_4_37 ( .A(sll_14_ML_int_4__37_), .B(sll_14_ML_int_4__21_), 
        .S(n204), .Z(sll_14_ML_int_5__37_) );
  MUX2_X1 sll_14_M1_4_38 ( .A(sll_14_ML_int_4__38_), .B(sll_14_ML_int_4__22_), 
        .S(n204), .Z(sll_14_ML_int_5__38_) );
  MUX2_X1 sll_14_M1_4_39 ( .A(sll_14_ML_int_4__39_), .B(sll_14_ML_int_4__23_), 
        .S(n204), .Z(sll_14_ML_int_5__39_) );
  MUX2_X1 sll_14_M1_4_40 ( .A(sll_14_ML_int_4__40_), .B(sll_14_ML_int_4__24_), 
        .S(n206), .Z(sll_14_ML_int_5__40_) );
  MUX2_X1 sll_14_M1_4_41 ( .A(sll_14_ML_int_4__41_), .B(sll_14_ML_int_4__25_), 
        .S(n206), .Z(sll_14_ML_int_5__41_) );
  MUX2_X1 sll_14_M1_4_42 ( .A(sll_14_ML_int_4__42_), .B(sll_14_ML_int_4__26_), 
        .S(n206), .Z(sll_14_ML_int_5__42_) );
  MUX2_X1 sll_14_M1_4_43 ( .A(sll_14_ML_int_4__43_), .B(sll_14_ML_int_4__27_), 
        .S(n206), .Z(sll_14_ML_int_5__43_) );
  MUX2_X1 sll_14_M1_4_44 ( .A(sll_14_ML_int_4__44_), .B(sll_14_ML_int_4__28_), 
        .S(n206), .Z(sll_14_ML_int_5__44_) );
  MUX2_X1 sll_14_M1_4_45 ( .A(sll_14_ML_int_4__45_), .B(sll_14_ML_int_4__29_), 
        .S(n206), .Z(sll_14_ML_int_5__45_) );
  MUX2_X1 sll_14_M1_4_46 ( .A(n220), .B(sll_14_ML_int_4__30_), .S(n206), .Z(
        sll_14_ML_int_5__46_) );
  MUX2_X1 sll_14_M1_5_32 ( .A(sll_14_ML_int_5__32_), .B(n248), .S(n199), .Z(
        N38) );
  MUX2_X1 sll_14_M1_5_33 ( .A(sll_14_ML_int_5__33_), .B(n241), .S(n200), .Z(
        N39) );
  MUX2_X1 sll_14_M1_5_34 ( .A(sll_14_ML_int_5__34_), .B(n3), .S(n199), .Z(N40)
         );
  MUX2_X1 sll_14_M1_5_35 ( .A(sll_14_ML_int_5__35_), .B(n2), .S(n199), .Z(N41)
         );
  MUX2_X1 sll_14_M1_5_36 ( .A(sll_14_ML_int_5__36_), .B(n246), .S(n200), .Z(
        N42) );
  MUX2_X1 sll_14_M1_5_37 ( .A(sll_14_ML_int_5__37_), .B(n239), .S(n200), .Z(
        N43) );
  MUX2_X1 sll_14_M1_5_38 ( .A(sll_14_ML_int_5__38_), .B(n243), .S(n200), .Z(
        N44) );
  MUX2_X1 sll_14_M1_5_39 ( .A(sll_14_ML_int_5__39_), .B(n236), .S(n199), .Z(
        N45) );
  MUX2_X1 sll_14_M1_5_40 ( .A(sll_14_ML_int_5__40_), .B(n247), .S(n199), .Z(
        N46) );
  MUX2_X1 sll_14_M1_5_41 ( .A(sll_14_ML_int_5__41_), .B(n240), .S(n200), .Z(
        N47) );
  MUX2_X1 sll_14_M1_5_42 ( .A(sll_14_ML_int_5__42_), .B(n244), .S(n200), .Z(
        N48) );
  MUX2_X1 sll_14_M1_5_43 ( .A(sll_14_ML_int_5__43_), .B(n237), .S(n200), .Z(
        N49) );
  MUX2_X1 sll_14_M1_5_44 ( .A(sll_14_ML_int_5__44_), .B(n245), .S(n200), .Z(
        N50) );
  MUX2_X1 sll_14_M1_5_45 ( .A(sll_14_ML_int_5__45_), .B(n238), .S(n200), .Z(
        N51) );
  MUX2_X1 sll_14_M1_5_46 ( .A(sll_14_ML_int_5__46_), .B(n242), .S(n199), .Z(
        N52) );
  MUX2_X1 sll_14_M1_5_47 ( .A(sll_14_ML_int_5__47_), .B(n235), .S(n199), .Z(
        N53) );
  MUX2_X1 sll_14_M1_5_48 ( .A(sll_14_ML_int_5__48_), .B(sll_14_ML_int_5__16_), 
        .S(n199), .Z(N54) );
  MUX2_X1 sll_14_M1_5_49 ( .A(sll_14_ML_int_5__49_), .B(sll_14_ML_int_5__17_), 
        .S(n199), .Z(N55) );
  MUX2_X1 sll_14_M1_5_50 ( .A(sll_14_ML_int_5__50_), .B(sll_14_ML_int_5__18_), 
        .S(n200), .Z(N56) );
  MUX2_X1 sll_14_M1_5_51 ( .A(sll_14_ML_int_5__51_), .B(sll_14_ML_int_5__19_), 
        .S(n199), .Z(N57) );
  MUX2_X1 sll_14_M1_5_52 ( .A(sll_14_ML_int_5__52_), .B(sll_14_ML_int_5__20_), 
        .S(n200), .Z(N58) );
  MUX2_X1 sll_14_M1_5_53 ( .A(sll_14_ML_int_5__53_), .B(sll_14_ML_int_5__21_), 
        .S(n199), .Z(N59) );
  MUX2_X1 sll_14_M1_5_54 ( .A(sll_14_ML_int_5__54_), .B(sll_14_ML_int_5__22_), 
        .S(n200), .Z(N60) );
  MUX2_X1 sll_14_M1_5_55 ( .A(sll_14_ML_int_5__55_), .B(sll_14_ML_int_5__23_), 
        .S(n199), .Z(N61) );
  MUX2_X1 sll_14_M1_5_56 ( .A(sll_14_ML_int_5__56_), .B(sll_14_ML_int_5__24_), 
        .S(n199), .Z(N62) );
  MUX2_X1 sll_14_M1_5_57 ( .A(sll_14_ML_int_5__57_), .B(sll_14_ML_int_5__25_), 
        .S(n199), .Z(N63) );
  MUX2_X1 sll_14_M1_5_58 ( .A(sll_14_ML_int_5__58_), .B(sll_14_ML_int_5__26_), 
        .S(n200), .Z(N64) );
  MUX2_X1 sll_14_M1_5_59 ( .A(sll_14_ML_int_5__59_), .B(sll_14_ML_int_5__27_), 
        .S(n200), .Z(N65) );
  MUX2_X1 sll_14_M1_5_60 ( .A(sll_14_ML_int_5__60_), .B(sll_14_ML_int_5__28_), 
        .S(n199), .Z(N66) );
  MUX2_X1 sll_14_M1_5_61 ( .A(sll_14_ML_int_5__61_), .B(sll_14_ML_int_5__29_), 
        .S(n200), .Z(N67) );
  MUX2_X1 sll_14_M1_5_62 ( .A(n220), .B(sll_14_ML_int_5__30_), .S(n200), .Z(
        N68) );
  DFF_X1 A_reg_63_ ( .D(n261), .CK(clk), .Q(result[63]) );
  XNOR2_X1 U3 ( .A(n32), .B(n165), .ZN(n_0_net__19_) );
  INV_X1 U4 ( .A(n202), .ZN(n201) );
  CLKBUF_X3 U5 ( .A(n217), .Z(n12) );
  INV_X1 U6 ( .A(N5), .ZN(n207) );
  INV_X1 U7 ( .A(n207), .ZN(n205) );
  INV_X2 U8 ( .A(n20), .ZN(n204) );
  BUF_X2 U9 ( .A(n181), .Z(n1) );
  INV_X1 U10 ( .A(n211), .ZN(n209) );
  AND2_X1 U11 ( .A1(sll_14_ML_int_4__3_), .A2(n207), .ZN(n2) );
  AND2_X1 U12 ( .A1(sll_14_ML_int_4__2_), .A2(n207), .ZN(n3) );
  XOR2_X1 U13 ( .A(N56), .B(n159), .Z(n_0_net__50_) );
  XOR2_X1 U14 ( .A(N61), .B(n164), .Z(n_0_net__55_) );
  XOR2_X1 U15 ( .A(N50), .B(n150), .Z(n_0_net__44_) );
  XOR2_X1 U16 ( .A(N54), .B(n157), .Z(n_0_net__48_) );
  XOR2_X1 U17 ( .A(N32), .B(n174), .Z(n_0_net__26_) );
  XOR2_X1 U18 ( .A(N48), .B(n148), .Z(n_0_net__42_) );
  AND3_X1 U19 ( .A1(N1), .A2(n67), .A3(N2), .ZN(n4) );
  AND3_X1 U20 ( .A1(N1), .A2(n67), .A3(N2), .ZN(n136) );
  CLKBUF_X1 U21 ( .A(n136), .Z(n5) );
  BUF_X1 U22 ( .A(sll_14_ML_int_1__2_), .Z(n11) );
  BUF_X1 U23 ( .A(sll_14_ML_int_2__1_), .Z(n6) );
  NOR2_X1 U24 ( .A1(n7), .A2(n8), .ZN(n15) );
  NAND2_X1 U25 ( .A1(n181), .A2(n180), .ZN(n7) );
  NAND2_X1 U26 ( .A1(n177), .A2(n176), .ZN(n8) );
  MUX2_X1 U27 ( .A(n17), .B(n11), .S(n1), .Z(n9) );
  BUF_X1 U28 ( .A(sll_14_ML_int_1__0_), .Z(n17) );
  CLKBUF_X1 U29 ( .A(n176), .Z(n13) );
  AND4_X1 U30 ( .A1(n5), .A2(N3), .A3(N5), .A4(n178), .ZN(n137) );
  BUF_X1 U31 ( .A(n177), .Z(n10) );
  INV_X2 U32 ( .A(n1), .ZN(n215) );
  BUF_X1 U33 ( .A(n180), .Z(n14) );
  NAND2_X1 U34 ( .A1(n15), .A2(sll_14_ML_int_1__0_), .ZN(n221) );
  AND2_X1 U35 ( .A1(sll_14_ML_int_4__3_), .A2(n16), .ZN(N9) );
  NOR2_X1 U36 ( .A1(n179), .A2(n201), .ZN(n16) );
  INV_X1 U37 ( .A(n182), .ZN(n217) );
  CLKBUF_X1 U38 ( .A(n212), .Z(n18) );
  AND2_X1 U39 ( .A1(n26), .A2(n14), .ZN(n19) );
  INV_X1 U40 ( .A(n205), .ZN(n20) );
  NAND4_X1 U41 ( .A1(n4), .A2(N3), .A3(N5), .A4(n178), .ZN(n21) );
  MUX2_X1 U42 ( .A(a[1]), .B(a[2]), .S(n182), .Z(sll_14_ML_int_1__2_) );
  AND2_X1 U43 ( .A1(sll_14_ML_int_2__0_), .A2(n14), .ZN(n22) );
  INV_X1 U44 ( .A(n66), .ZN(n23) );
  AND2_X1 U45 ( .A1(sll_14_ML_int_4__2_), .A2(n24), .ZN(N8) );
  AND2_X1 U46 ( .A1(n13), .A2(n25), .ZN(n24) );
  INV_X1 U47 ( .A(i_5_), .ZN(n25) );
  NAND2_X1 U48 ( .A1(n19), .A2(sll_14_ML_int_2__1_), .ZN(n228) );
  AND2_X1 U49 ( .A1(n211), .A2(n208), .ZN(n26) );
  XNOR2_X1 U50 ( .A(n27), .B(n146), .ZN(n_0_net__4_) );
  OR2_X1 U51 ( .A1(n199), .A2(n229), .ZN(n27) );
  XNOR2_X1 U52 ( .A(N6), .B(n21), .ZN(n_0_net__0_) );
  INV_X1 U53 ( .A(n221), .ZN(n248) );
  BUF_X1 U54 ( .A(n191), .Z(n195) );
  BUF_X1 U55 ( .A(n191), .Z(n194) );
  BUF_X1 U56 ( .A(n191), .Z(n193) );
  BUF_X1 U57 ( .A(n192), .Z(n197) );
  BUF_X1 U58 ( .A(n192), .Z(n196) );
  BUF_X1 U59 ( .A(n183), .Z(n186) );
  BUF_X1 U60 ( .A(n183), .Z(n187) );
  BUF_X1 U61 ( .A(n184), .Z(n188) );
  BUF_X1 U62 ( .A(n184), .Z(n189) );
  BUF_X1 U63 ( .A(n183), .Z(n185) );
  XNOR2_X1 U64 ( .A(n28), .B(n151), .ZN(n_0_net__13_) );
  OR2_X1 U65 ( .A1(n200), .A2(n225), .ZN(n28) );
  XNOR2_X1 U66 ( .A(N40), .B(n169), .ZN(n_0_net__34_) );
  XNOR2_X1 U67 ( .A(N38), .B(n169), .ZN(n_0_net__32_) );
  INV_X1 U68 ( .A(n222), .ZN(n244) );
  INV_X1 U69 ( .A(n229), .ZN(n246) );
  INV_X1 U70 ( .A(n223), .ZN(n237) );
  INV_X1 U71 ( .A(n224), .ZN(n245) );
  INV_X1 U72 ( .A(n233), .ZN(n247) );
  INV_X1 U73 ( .A(n225), .ZN(n238) );
  INV_X1 U74 ( .A(n234), .ZN(n240) );
  INV_X1 U75 ( .A(n230), .ZN(n239) );
  INV_X1 U76 ( .A(n231), .ZN(n243) );
  INV_X1 U77 ( .A(n232), .ZN(n236) );
  CLKBUF_X1 U78 ( .A(n66), .Z(n68) );
  CLKBUF_X1 U79 ( .A(n12), .Z(n66) );
  NOR2_X1 U80 ( .A1(n325), .A2(n190), .ZN(n70) );
  MUX2_X1 U81 ( .A(sll_14_ML_int_2__0_), .B(sll_14_ML_int_2__4_), .S(n214), 
        .Z(sll_14_ML_int_3__4_) );
  MUX2_X1 U82 ( .A(n17), .B(sll_14_ML_int_1__2_), .S(n1), .Z(
        sll_14_ML_int_2__2_) );
  INV_X1 U83 ( .A(n202), .ZN(n199) );
  INV_X1 U84 ( .A(n20), .ZN(n206) );
  XNOR2_X1 U85 ( .A(n29), .B(n170), .ZN(n_0_net__22_) );
  NAND2_X1 U86 ( .A1(sll_14_ML_int_5__22_), .A2(n203), .ZN(n29) );
  XNOR2_X1 U87 ( .A(n30), .B(n167), .ZN(n_0_net__21_) );
  NAND2_X1 U88 ( .A1(sll_14_ML_int_5__21_), .A2(n203), .ZN(n30) );
  XNOR2_X1 U89 ( .A(n31), .B(n166), .ZN(n_0_net__20_) );
  NAND2_X1 U90 ( .A1(sll_14_ML_int_5__20_), .A2(n203), .ZN(n31) );
  NAND2_X1 U91 ( .A1(sll_14_ML_int_5__19_), .A2(n203), .ZN(n32) );
  INV_X1 U92 ( .A(n211), .ZN(n210) );
  MUX2_X1 U93 ( .A(sll_14_ML_int_1__1_), .B(sll_14_ML_int_1__3_), .S(n1), .Z(
        sll_14_ML_int_2__3_) );
  XNOR2_X1 U94 ( .A(n33), .B(n162), .ZN(n_0_net__16_) );
  NAND2_X1 U95 ( .A1(sll_14_ML_int_5__16_), .A2(n203), .ZN(n33) );
  XNOR2_X1 U96 ( .A(n34), .B(n163), .ZN(n_0_net__17_) );
  NAND2_X1 U97 ( .A1(sll_14_ML_int_5__17_), .A2(n203), .ZN(n34) );
  XNOR2_X1 U98 ( .A(n35), .B(n164), .ZN(n_0_net__18_) );
  NAND2_X1 U99 ( .A1(sll_14_ML_int_5__18_), .A2(n203), .ZN(n35) );
  INV_X1 U100 ( .A(n226), .ZN(n242) );
  INV_X1 U101 ( .A(n227), .ZN(n235) );
  INV_X1 U102 ( .A(n202), .ZN(n200) );
  NOR2_X1 U103 ( .A1(N74), .A2(n325), .ZN(n71) );
  INV_X1 U104 ( .A(n135), .ZN(n325) );
  AND2_X1 U105 ( .A1(N76), .A2(n135), .ZN(N147) );
  AND2_X1 U106 ( .A1(N77), .A2(n135), .ZN(N148) );
  AND2_X1 U107 ( .A1(N78), .A2(n135), .ZN(N149) );
  AND2_X1 U108 ( .A1(N79), .A2(n135), .ZN(N150) );
  AND2_X1 U109 ( .A1(N80), .A2(n135), .ZN(N151) );
  INV_X1 U110 ( .A(n72), .ZN(n262) );
  AOI22_X1 U111 ( .A1(tempResult[62]), .A2(n198), .B1(result[62]), .B2(n185), 
        .ZN(n72) );
  INV_X1 U112 ( .A(n73), .ZN(n263) );
  AOI22_X1 U113 ( .A1(tempResult[61]), .A2(n198), .B1(result[61]), .B2(n185), 
        .ZN(n73) );
  INV_X1 U114 ( .A(n74), .ZN(n264) );
  AOI22_X1 U115 ( .A1(tempResult[60]), .A2(n198), .B1(result[60]), .B2(n185), 
        .ZN(n74) );
  INV_X1 U116 ( .A(n83), .ZN(n273) );
  AOI22_X1 U117 ( .A1(tempResult[51]), .A2(n197), .B1(result[51]), .B2(n186), 
        .ZN(n83) );
  INV_X1 U118 ( .A(n85), .ZN(n275) );
  AOI22_X1 U119 ( .A1(tempResult[49]), .A2(n197), .B1(result[49]), .B2(n186), 
        .ZN(n85) );
  BUF_X1 U120 ( .A(a[31]), .Z(n218) );
  INV_X1 U121 ( .A(N5), .ZN(n208) );
  INV_X1 U122 ( .A(n84), .ZN(n274) );
  AOI22_X1 U123 ( .A1(tempResult[50]), .A2(n197), .B1(result[50]), .B2(n186), 
        .ZN(n84) );
  INV_X1 U124 ( .A(n75), .ZN(n265) );
  AOI22_X1 U125 ( .A1(tempResult[59]), .A2(n197), .B1(result[59]), .B2(n185), 
        .ZN(n75) );
  INV_X1 U126 ( .A(n76), .ZN(n266) );
  AOI22_X1 U127 ( .A1(tempResult[58]), .A2(n197), .B1(result[58]), .B2(n185), 
        .ZN(n76) );
  INV_X1 U128 ( .A(n77), .ZN(n267) );
  AOI22_X1 U129 ( .A1(tempResult[57]), .A2(n197), .B1(result[57]), .B2(n185), 
        .ZN(n77) );
  INV_X1 U130 ( .A(n78), .ZN(n268) );
  AOI22_X1 U131 ( .A1(tempResult[56]), .A2(n197), .B1(result[56]), .B2(n185), 
        .ZN(n78) );
  INV_X1 U132 ( .A(n79), .ZN(n269) );
  AOI22_X1 U133 ( .A1(tempResult[55]), .A2(n197), .B1(result[55]), .B2(n185), 
        .ZN(n79) );
  INV_X1 U134 ( .A(n80), .ZN(n270) );
  AOI22_X1 U135 ( .A1(tempResult[54]), .A2(n197), .B1(result[54]), .B2(n185), 
        .ZN(n80) );
  INV_X1 U136 ( .A(n81), .ZN(n271) );
  AOI22_X1 U137 ( .A1(tempResult[53]), .A2(n197), .B1(result[53]), .B2(n185), 
        .ZN(n81) );
  INV_X1 U138 ( .A(n86), .ZN(n276) );
  AOI22_X1 U139 ( .A1(tempResult[48]), .A2(n197), .B1(result[48]), .B2(n186), 
        .ZN(n86) );
  INV_X1 U140 ( .A(n87), .ZN(n277) );
  AOI22_X1 U141 ( .A1(tempResult[47]), .A2(n196), .B1(result[47]), .B2(n186), 
        .ZN(n87) );
  INV_X1 U142 ( .A(n88), .ZN(n278) );
  AOI22_X1 U143 ( .A1(tempResult[46]), .A2(n196), .B1(result[46]), .B2(n186), 
        .ZN(n88) );
  INV_X1 U157 ( .A(n82), .ZN(n272) );
  AOI22_X1 U162 ( .A1(tempResult[52]), .A2(n197), .B1(result[52]), .B2(n185), 
        .ZN(n82) );
  INV_X1 U163 ( .A(n89), .ZN(n279) );
  AOI22_X1 U165 ( .A1(tempResult[45]), .A2(n196), .B1(result[45]), .B2(n186), 
        .ZN(n89) );
  INV_X1 U169 ( .A(n90), .ZN(n280) );
  AOI22_X1 U171 ( .A1(tempResult[44]), .A2(n196), .B1(result[44]), .B2(n186), 
        .ZN(n90) );
  INV_X1 U180 ( .A(n91), .ZN(n281) );
  AOI22_X1 U182 ( .A1(tempResult[43]), .A2(n196), .B1(result[43]), .B2(n186), 
        .ZN(n91) );
  INV_X1 U189 ( .A(n92), .ZN(n282) );
  AOI22_X1 U193 ( .A1(tempResult[42]), .A2(n196), .B1(result[42]), .B2(n186), 
        .ZN(n92) );
  INV_X1 U194 ( .A(n93), .ZN(n283) );
  AOI22_X1 U195 ( .A1(tempResult[41]), .A2(n196), .B1(result[41]), .B2(n186), 
        .ZN(n93) );
  INV_X1 U197 ( .A(n94), .ZN(n284) );
  AOI22_X1 U198 ( .A1(tempResult[40]), .A2(n196), .B1(result[40]), .B2(n186), 
        .ZN(n94) );
  INV_X1 U199 ( .A(n95), .ZN(n285) );
  AOI22_X1 U200 ( .A1(tempResult[39]), .A2(n196), .B1(result[39]), .B2(n187), 
        .ZN(n95) );
  INV_X1 U203 ( .A(n96), .ZN(n286) );
  AOI22_X1 U207 ( .A1(tempResult[38]), .A2(n196), .B1(result[38]), .B2(n187), 
        .ZN(n96) );
  INV_X1 U208 ( .A(n97), .ZN(n287) );
  AOI22_X1 U209 ( .A1(tempResult[37]), .A2(n196), .B1(result[37]), .B2(n187), 
        .ZN(n97) );
  INV_X1 U210 ( .A(n98), .ZN(n288) );
  AOI22_X1 U211 ( .A1(tempResult[36]), .A2(n196), .B1(result[36]), .B2(n187), 
        .ZN(n98) );
  INV_X1 U212 ( .A(n99), .ZN(n289) );
  AOI22_X1 U213 ( .A1(tempResult[35]), .A2(n195), .B1(result[35]), .B2(n187), 
        .ZN(n99) );
  INV_X1 U214 ( .A(n114), .ZN(n304) );
  AOI22_X1 U215 ( .A1(tempResult[20]), .A2(n194), .B1(result[20]), .B2(n188), 
        .ZN(n114) );
  BUF_X1 U216 ( .A(a[31]), .Z(n219) );
  BUF_X1 U217 ( .A(a[31]), .Z(n220) );
  INV_X1 U218 ( .A(n101), .ZN(n291) );
  AOI22_X1 U219 ( .A1(tempResult[33]), .A2(n195), .B1(result[33]), .B2(n187), 
        .ZN(n101) );
  INV_X1 U220 ( .A(n111), .ZN(n301) );
  AOI22_X1 U221 ( .A1(tempResult[23]), .A2(n194), .B1(result[23]), .B2(n188), 
        .ZN(n111) );
  INV_X1 U222 ( .A(n100), .ZN(n290) );
  AOI22_X1 U223 ( .A1(tempResult[34]), .A2(n195), .B1(result[34]), .B2(n187), 
        .ZN(n100) );
  INV_X1 U224 ( .A(n102), .ZN(n292) );
  AOI22_X1 U225 ( .A1(tempResult[32]), .A2(n195), .B1(result[32]), .B2(n187), 
        .ZN(n102) );
  INV_X1 U226 ( .A(n103), .ZN(n293) );
  AOI22_X1 U227 ( .A1(tempResult[31]), .A2(n195), .B1(result[31]), .B2(n187), 
        .ZN(n103) );
  INV_X1 U228 ( .A(n104), .ZN(n294) );
  AOI22_X1 U229 ( .A1(tempResult[30]), .A2(n195), .B1(result[30]), .B2(n187), 
        .ZN(n104) );
  INV_X1 U230 ( .A(n105), .ZN(n295) );
  AOI22_X1 U231 ( .A1(tempResult[29]), .A2(n195), .B1(result[29]), .B2(n187), 
        .ZN(n105) );
  INV_X1 U232 ( .A(n106), .ZN(n296) );
  AOI22_X1 U233 ( .A1(tempResult[28]), .A2(n195), .B1(result[28]), .B2(n187), 
        .ZN(n106) );
  INV_X1 U234 ( .A(n107), .ZN(n297) );
  AOI22_X1 U235 ( .A1(tempResult[27]), .A2(n195), .B1(result[27]), .B2(n188), 
        .ZN(n107) );
  INV_X1 U236 ( .A(n108), .ZN(n298) );
  AOI22_X1 U237 ( .A1(tempResult[26]), .A2(n195), .B1(result[26]), .B2(n188), 
        .ZN(n108) );
  INV_X1 U238 ( .A(n109), .ZN(n299) );
  AOI22_X1 U239 ( .A1(tempResult[25]), .A2(n195), .B1(result[25]), .B2(n188), 
        .ZN(n109) );
  INV_X1 U240 ( .A(n110), .ZN(n300) );
  AOI22_X1 U241 ( .A1(tempResult[24]), .A2(n195), .B1(result[24]), .B2(n188), 
        .ZN(n110) );
  INV_X1 U242 ( .A(n112), .ZN(n302) );
  AOI22_X1 U243 ( .A1(tempResult[22]), .A2(n194), .B1(result[22]), .B2(n188), 
        .ZN(n112) );
  INV_X1 U244 ( .A(n113), .ZN(n303) );
  AOI22_X1 U245 ( .A1(tempResult[21]), .A2(n194), .B1(result[21]), .B2(n188), 
        .ZN(n113) );
  INV_X1 U246 ( .A(n121), .ZN(n311) );
  AOI22_X1 U247 ( .A1(tempResult[13]), .A2(n194), .B1(result[13]), .B2(n189), 
        .ZN(n121) );
  INV_X1 U248 ( .A(n131), .ZN(n321) );
  AOI22_X1 U249 ( .A1(tempResult[3]), .A2(n193), .B1(result[3]), .B2(n190), 
        .ZN(n131) );
  INV_X1 U250 ( .A(n132), .ZN(n322) );
  AOI22_X1 U251 ( .A1(tempResult[2]), .A2(n193), .B1(result[2]), .B2(n190), 
        .ZN(n132) );
  INV_X1 U252 ( .A(n133), .ZN(n323) );
  AOI22_X1 U253 ( .A1(tempResult[1]), .A2(n193), .B1(result[1]), .B2(n190), 
        .ZN(n133) );
  INV_X1 U254 ( .A(n134), .ZN(n324) );
  AOI22_X1 U255 ( .A1(tempResult[0]), .A2(n193), .B1(result[0]), .B2(n190), 
        .ZN(n134) );
  INV_X1 U256 ( .A(n116), .ZN(n306) );
  AOI22_X1 U257 ( .A1(tempResult[18]), .A2(n194), .B1(result[18]), .B2(n188), 
        .ZN(n116) );
  INV_X1 U258 ( .A(n117), .ZN(n307) );
  AOI22_X1 U259 ( .A1(tempResult[17]), .A2(n194), .B1(result[17]), .B2(n188), 
        .ZN(n117) );
  INV_X1 U260 ( .A(n118), .ZN(n308) );
  AOI22_X1 U261 ( .A1(tempResult[16]), .A2(n194), .B1(result[16]), .B2(n188), 
        .ZN(n118) );
  INV_X1 U262 ( .A(n119), .ZN(n309) );
  AOI22_X1 U263 ( .A1(tempResult[15]), .A2(n194), .B1(result[15]), .B2(n189), 
        .ZN(n119) );
  INV_X1 U264 ( .A(n123), .ZN(n313) );
  AOI22_X1 U265 ( .A1(tempResult[11]), .A2(n193), .B1(result[11]), .B2(n189), 
        .ZN(n123) );
  INV_X1 U266 ( .A(n124), .ZN(n314) );
  AOI22_X1 U267 ( .A1(tempResult[10]), .A2(n193), .B1(result[10]), .B2(n189), 
        .ZN(n124) );
  INV_X1 U268 ( .A(n125), .ZN(n315) );
  AOI22_X1 U269 ( .A1(tempResult[9]), .A2(n193), .B1(result[9]), .B2(n189), 
        .ZN(n125) );
  INV_X1 U270 ( .A(n126), .ZN(n316) );
  AOI22_X1 U271 ( .A1(tempResult[8]), .A2(n193), .B1(result[8]), .B2(n189), 
        .ZN(n126) );
  INV_X1 U272 ( .A(n127), .ZN(n317) );
  AOI22_X1 U273 ( .A1(tempResult[7]), .A2(n193), .B1(result[7]), .B2(n189), 
        .ZN(n127) );
  INV_X1 U274 ( .A(n115), .ZN(n305) );
  AOI22_X1 U275 ( .A1(tempResult[19]), .A2(n194), .B1(result[19]), .B2(n188), 
        .ZN(n115) );
  INV_X1 U276 ( .A(n120), .ZN(n310) );
  AOI22_X1 U277 ( .A1(tempResult[14]), .A2(n194), .B1(result[14]), .B2(n189), 
        .ZN(n120) );
  INV_X1 U278 ( .A(n122), .ZN(n312) );
  AOI22_X1 U279 ( .A1(tempResult[12]), .A2(n194), .B1(result[12]), .B2(n189), 
        .ZN(n122) );
  INV_X1 U280 ( .A(n128), .ZN(n318) );
  AOI22_X1 U281 ( .A1(tempResult[6]), .A2(n193), .B1(result[6]), .B2(n189), 
        .ZN(n128) );
  INV_X1 U282 ( .A(n129), .ZN(n319) );
  AOI22_X1 U283 ( .A1(tempResult[5]), .A2(n193), .B1(result[5]), .B2(n189), 
        .ZN(n129) );
  INV_X1 U284 ( .A(n130), .ZN(n320) );
  AOI22_X1 U285 ( .A1(tempResult[4]), .A2(n193), .B1(result[4]), .B2(n189), 
        .ZN(n130) );
  NOR2_X1 U286 ( .A1(reset), .A2(n200), .ZN(n135) );
  MUX2_X1 U287 ( .A(b[30]), .B(b[31]), .S(n68), .Z(n36) );
  MUX2_X1 U288 ( .A(b[28]), .B(b[29]), .S(n68), .Z(n37) );
  MUX2_X1 U289 ( .A(n37), .B(n36), .S(n216), .Z(n38) );
  MUX2_X1 U290 ( .A(b[26]), .B(b[27]), .S(n68), .Z(n39) );
  MUX2_X1 U291 ( .A(b[24]), .B(b[25]), .S(n68), .Z(n40) );
  MUX2_X1 U292 ( .A(n40), .B(n39), .S(n216), .Z(n41) );
  MUX2_X1 U293 ( .A(n41), .B(n38), .S(n213), .Z(n42) );
  MUX2_X1 U294 ( .A(b[22]), .B(b[23]), .S(n68), .Z(n43) );
  MUX2_X1 U295 ( .A(b[20]), .B(b[21]), .S(n68), .Z(n44) );
  MUX2_X1 U296 ( .A(n44), .B(n43), .S(n216), .Z(n45) );
  MUX2_X1 U297 ( .A(b[18]), .B(b[19]), .S(n68), .Z(n46) );
  MUX2_X1 U298 ( .A(b[16]), .B(b[17]), .S(n68), .Z(n47) );
  MUX2_X1 U299 ( .A(n47), .B(n46), .S(n216), .Z(n48) );
  MUX2_X1 U300 ( .A(n48), .B(n45), .S(n213), .Z(n49) );
  MUX2_X1 U301 ( .A(n49), .B(n42), .S(n210), .Z(n50) );
  MUX2_X1 U302 ( .A(b[14]), .B(b[15]), .S(n68), .Z(n51) );
  MUX2_X1 U303 ( .A(b[12]), .B(b[13]), .S(n68), .Z(n52) );
  MUX2_X1 U304 ( .A(n52), .B(n51), .S(n216), .Z(n53) );
  MUX2_X1 U305 ( .A(b[10]), .B(b[11]), .S(n68), .Z(n54) );
  MUX2_X1 U306 ( .A(b[8]), .B(b[9]), .S(n68), .Z(n55) );
  MUX2_X1 U307 ( .A(n55), .B(n54), .S(n216), .Z(n56) );
  MUX2_X1 U308 ( .A(n56), .B(n53), .S(n213), .Z(n57) );
  MUX2_X1 U309 ( .A(b[6]), .B(b[7]), .S(n66), .Z(n58) );
  MUX2_X1 U310 ( .A(b[4]), .B(b[5]), .S(n66), .Z(n59) );
  MUX2_X1 U311 ( .A(n59), .B(n58), .S(n216), .Z(n60) );
  MUX2_X1 U312 ( .A(b[2]), .B(b[3]), .S(n66), .Z(n61) );
  MUX2_X1 U313 ( .A(b[0]), .B(b[1]), .S(n66), .Z(n62) );
  MUX2_X1 U314 ( .A(n62), .B(n61), .S(n216), .Z(n63) );
  MUX2_X1 U315 ( .A(n63), .B(n60), .S(n213), .Z(n64) );
  MUX2_X1 U316 ( .A(n64), .B(n57), .S(n210), .Z(n65) );
  MUX2_X1 U317 ( .A(n65), .B(n50), .S(n204), .Z(N74) );
  CLKBUF_X1 U318 ( .A(n137), .Z(n138) );
  CLKBUF_X1 U319 ( .A(n137), .Z(n139) );
  INV_X1 U320 ( .A(n137), .ZN(n140) );
  INV_X1 U321 ( .A(n137), .ZN(n141) );
  INV_X1 U322 ( .A(n140), .ZN(n142) );
  INV_X1 U323 ( .A(n140), .ZN(n143) );
  INV_X1 U324 ( .A(n141), .ZN(n144) );
  INV_X1 U325 ( .A(n140), .ZN(n145) );
  INV_X1 U326 ( .A(n141), .ZN(n146) );
  INV_X1 U327 ( .A(n140), .ZN(n147) );
  INV_X1 U328 ( .A(n141), .ZN(n148) );
  INV_X1 U329 ( .A(n140), .ZN(n149) );
  INV_X1 U330 ( .A(n141), .ZN(n150) );
  INV_X1 U331 ( .A(n141), .ZN(n151) );
  INV_X1 U332 ( .A(n140), .ZN(n152) );
  INV_X1 U333 ( .A(n138), .ZN(n153) );
  INV_X1 U334 ( .A(n138), .ZN(n154) );
  INV_X1 U335 ( .A(n138), .ZN(n155) );
  INV_X1 U336 ( .A(n153), .ZN(n156) );
  INV_X1 U337 ( .A(n153), .ZN(n157) );
  INV_X1 U338 ( .A(n153), .ZN(n158) );
  INV_X1 U339 ( .A(n153), .ZN(n159) );
  INV_X1 U340 ( .A(n154), .ZN(n160) );
  INV_X1 U341 ( .A(n154), .ZN(n161) );
  INV_X1 U342 ( .A(n154), .ZN(n162) );
  INV_X1 U343 ( .A(n154), .ZN(n163) );
  INV_X1 U344 ( .A(n155), .ZN(n164) );
  INV_X1 U345 ( .A(n155), .ZN(n165) );
  INV_X1 U346 ( .A(n155), .ZN(n166) );
  INV_X1 U347 ( .A(n155), .ZN(n167) );
  INV_X1 U348 ( .A(n139), .ZN(n168) );
  INV_X1 U349 ( .A(n139), .ZN(n169) );
  INV_X1 U350 ( .A(n168), .ZN(n170) );
  INV_X1 U351 ( .A(n168), .ZN(n171) );
  INV_X1 U352 ( .A(n168), .ZN(n172) );
  INV_X1 U353 ( .A(n168), .ZN(n173) );
  INV_X1 U354 ( .A(n168), .ZN(n174) );
  INV_X1 U355 ( .A(n169), .ZN(n175) );
  INV_X1 U356 ( .A(n228), .ZN(n241) );
  INV_X1 U357 ( .A(n10), .ZN(n178) );
  INV_X1 U358 ( .A(n13), .ZN(n179) );
  INV_X1 U359 ( .A(N3), .ZN(n214) );
  INV_X1 U360 ( .A(n1), .ZN(n216) );
  AOI22_X1 U361 ( .A1(tempResult[63]), .A2(n198), .B1(result[63]), .B2(n185), 
        .ZN(n69) );
  AND2_X1 U362 ( .A1(n23), .A2(n135), .ZN(N146) );
  INV_X1 U363 ( .A(n69), .ZN(n261) );
  BUF_X1 U364 ( .A(n71), .Z(n183) );
  BUF_X1 U365 ( .A(n71), .Z(n184) );
  BUF_X1 U366 ( .A(n184), .Z(n190) );
  BUF_X1 U367 ( .A(n70), .Z(n191) );
  BUF_X1 U368 ( .A(n70), .Z(n192) );
  BUF_X1 U369 ( .A(n192), .Z(n198) );
  INV_X1 U370 ( .A(i_5_), .ZN(n202) );
  INV_X1 U371 ( .A(i_5_), .ZN(n203) );
  INV_X1 U372 ( .A(N4), .ZN(n211) );
  INV_X1 U373 ( .A(N4), .ZN(n212) );
  INV_X4 U374 ( .A(n214), .ZN(n213) );
  AND2_X1 U375 ( .A1(n182), .A2(a[0]), .ZN(sll_14_ML_int_1__0_) );
  AND2_X1 U376 ( .A1(sll_14_ML_int_1__0_), .A2(n1), .ZN(sll_14_ML_int_2__0_)
         );
  AND2_X1 U377 ( .A1(sll_14_ML_int_1__1_), .A2(n1), .ZN(sll_14_ML_int_2__1_)
         );
  AND2_X1 U378 ( .A1(n6), .A2(n14), .ZN(sll_14_ML_int_3__1_) );
  AND2_X1 U379 ( .A1(sll_14_ML_int_2__2_), .A2(n214), .ZN(sll_14_ML_int_3__2_)
         );
  AND2_X1 U380 ( .A1(sll_14_ML_int_2__3_), .A2(n214), .ZN(sll_14_ML_int_3__3_)
         );
  AND2_X1 U381 ( .A1(n22), .A2(n18), .ZN(sll_14_ML_int_4__0_) );
  AND2_X1 U382 ( .A1(sll_14_ML_int_3__1_), .A2(n18), .ZN(sll_14_ML_int_4__1_)
         );
  AND2_X1 U383 ( .A1(sll_14_ML_int_3__2_), .A2(n18), .ZN(sll_14_ML_int_4__2_)
         );
  AND2_X1 U384 ( .A1(sll_14_ML_int_3__3_), .A2(n18), .ZN(sll_14_ML_int_4__3_)
         );
  AND2_X1 U385 ( .A1(sll_14_ML_int_3__4_), .A2(n212), .ZN(sll_14_ML_int_4__4_)
         );
  AND2_X1 U386 ( .A1(sll_14_ML_int_3__5_), .A2(n212), .ZN(sll_14_ML_int_4__5_)
         );
  AND2_X1 U387 ( .A1(sll_14_ML_int_3__6_), .A2(n212), .ZN(sll_14_ML_int_4__6_)
         );
  AND2_X1 U388 ( .A1(sll_14_ML_int_3__7_), .A2(n212), .ZN(sll_14_ML_int_4__7_)
         );
  NAND2_X1 U389 ( .A1(sll_14_ML_int_4__10_), .A2(n20), .ZN(n222) );
  NAND2_X1 U390 ( .A1(sll_14_ML_int_4__11_), .A2(n20), .ZN(n223) );
  NAND2_X1 U391 ( .A1(sll_14_ML_int_4__12_), .A2(n20), .ZN(n224) );
  NAND2_X1 U392 ( .A1(sll_14_ML_int_4__13_), .A2(n207), .ZN(n225) );
  NAND2_X1 U393 ( .A1(sll_14_ML_int_4__14_), .A2(n207), .ZN(n226) );
  NAND2_X1 U394 ( .A1(sll_14_ML_int_4__15_), .A2(n207), .ZN(n227) );
  NAND2_X1 U395 ( .A1(sll_14_ML_int_4__4_), .A2(n207), .ZN(n229) );
  NAND2_X1 U396 ( .A1(sll_14_ML_int_4__5_), .A2(n207), .ZN(n230) );
  NAND2_X1 U397 ( .A1(sll_14_ML_int_4__6_), .A2(n20), .ZN(n231) );
  NAND2_X1 U398 ( .A1(sll_14_ML_int_4__7_), .A2(n20), .ZN(n232) );
  NAND2_X1 U399 ( .A1(sll_14_ML_int_4__8_), .A2(n20), .ZN(n233) );
  NAND2_X1 U400 ( .A1(sll_14_ML_int_4__9_), .A2(n20), .ZN(n234) );
  NOR2_X1 U401 ( .A1(n221), .A2(i_5_), .ZN(N6) );
  NOR2_X1 U402 ( .A1(n199), .A2(n222), .ZN(N16) );
  NOR2_X1 U403 ( .A1(n200), .A2(n223), .ZN(N17) );
  NOR2_X1 U404 ( .A1(n199), .A2(n224), .ZN(N18) );
  NOR2_X1 U405 ( .A1(n199), .A2(n226), .ZN(N20) );
  NOR2_X1 U406 ( .A1(n200), .A2(n227), .ZN(N21) );
  NOR2_X1 U407 ( .A1(n201), .A2(n228), .ZN(N7) );
  AND2_X1 U408 ( .A1(sll_14_ML_int_5__23_), .A2(n203), .ZN(N29) );
  AND2_X1 U409 ( .A1(sll_14_ML_int_5__24_), .A2(n203), .ZN(N30) );
  AND2_X1 U410 ( .A1(sll_14_ML_int_5__25_), .A2(n203), .ZN(N31) );
  AND2_X1 U411 ( .A1(sll_14_ML_int_5__26_), .A2(n203), .ZN(N32) );
  AND2_X1 U412 ( .A1(sll_14_ML_int_5__27_), .A2(n203), .ZN(N33) );
  AND2_X1 U413 ( .A1(sll_14_ML_int_5__28_), .A2(n203), .ZN(N34) );
  AND2_X1 U414 ( .A1(sll_14_ML_int_5__29_), .A2(n203), .ZN(N35) );
  AND2_X1 U415 ( .A1(sll_14_ML_int_5__30_), .A2(n203), .ZN(N36) );
  AND2_X1 U416 ( .A1(sll_14_ML_int_5__31_), .A2(n203), .ZN(N37) );
  NOR2_X1 U417 ( .A1(n200), .A2(n230), .ZN(N11) );
  NOR2_X1 U418 ( .A1(n199), .A2(n231), .ZN(N12) );
  NOR2_X1 U419 ( .A1(n200), .A2(n232), .ZN(N13) );
  NOR2_X1 U420 ( .A1(n199), .A2(n233), .ZN(N14) );
  NOR2_X1 U421 ( .A1(n200), .A2(n234), .ZN(N15) );
  MUX2_X1 U422 ( .A(n220), .B(n249), .S(n206), .Z(sll_14_ML_int_5__47_) );
  MUX2_X1 U423 ( .A(n220), .B(sll_14_ML_int_4__32_), .S(n204), .Z(
        sll_14_ML_int_5__48_) );
  MUX2_X1 U424 ( .A(n250), .B(sll_14_ML_int_3__24_), .S(n209), .Z(
        sll_14_ML_int_4__32_) );
  MUX2_X1 U425 ( .A(n220), .B(sll_14_ML_int_4__33_), .S(n204), .Z(
        sll_14_ML_int_5__49_) );
  MUX2_X1 U426 ( .A(n251), .B(sll_14_ML_int_3__25_), .S(n209), .Z(
        sll_14_ML_int_4__33_) );
  MUX2_X1 U427 ( .A(n220), .B(sll_14_ML_int_4__34_), .S(n204), .Z(
        sll_14_ML_int_5__50_) );
  MUX2_X1 U428 ( .A(n252), .B(sll_14_ML_int_3__26_), .S(n209), .Z(
        sll_14_ML_int_4__34_) );
  MUX2_X1 U429 ( .A(n220), .B(sll_14_ML_int_4__35_), .S(n204), .Z(
        sll_14_ML_int_5__51_) );
  MUX2_X1 U430 ( .A(n253), .B(sll_14_ML_int_3__27_), .S(n209), .Z(
        sll_14_ML_int_4__35_) );
  MUX2_X1 U431 ( .A(n220), .B(sll_14_ML_int_4__36_), .S(n204), .Z(
        sll_14_ML_int_5__52_) );
  MUX2_X1 U432 ( .A(n254), .B(sll_14_ML_int_3__28_), .S(n210), .Z(
        sll_14_ML_int_4__36_) );
  MUX2_X1 U433 ( .A(n220), .B(sll_14_ML_int_4__37_), .S(n204), .Z(
        sll_14_ML_int_5__53_) );
  MUX2_X1 U434 ( .A(n255), .B(sll_14_ML_int_3__29_), .S(n210), .Z(
        sll_14_ML_int_4__37_) );
  MUX2_X1 U435 ( .A(n220), .B(sll_14_ML_int_4__38_), .S(n204), .Z(
        sll_14_ML_int_5__54_) );
  MUX2_X1 U436 ( .A(n220), .B(sll_14_ML_int_3__30_), .S(n209), .Z(
        sll_14_ML_int_4__38_) );
  MUX2_X1 U437 ( .A(n219), .B(sll_14_ML_int_4__39_), .S(n206), .Z(
        sll_14_ML_int_5__55_) );
  MUX2_X1 U438 ( .A(n219), .B(n256), .S(n210), .Z(sll_14_ML_int_4__39_) );
  MUX2_X1 U439 ( .A(n219), .B(sll_14_ML_int_4__40_), .S(n206), .Z(
        sll_14_ML_int_5__56_) );
  MUX2_X1 U440 ( .A(n219), .B(n250), .S(n210), .Z(sll_14_ML_int_4__40_) );
  MUX2_X1 U441 ( .A(n257), .B(sll_14_ML_int_2__28_), .S(n213), .Z(n250) );
  MUX2_X1 U442 ( .A(n219), .B(sll_14_ML_int_4__41_), .S(n206), .Z(
        sll_14_ML_int_5__57_) );
  MUX2_X1 U443 ( .A(n219), .B(n251), .S(n210), .Z(sll_14_ML_int_4__41_) );
  MUX2_X1 U444 ( .A(n258), .B(sll_14_ML_int_2__29_), .S(n213), .Z(n251) );
  MUX2_X1 U445 ( .A(n219), .B(sll_14_ML_int_4__42_), .S(n204), .Z(
        sll_14_ML_int_5__58_) );
  MUX2_X1 U446 ( .A(n219), .B(n252), .S(n210), .Z(sll_14_ML_int_4__42_) );
  MUX2_X1 U447 ( .A(n219), .B(sll_14_ML_int_2__30_), .S(n213), .Z(n252) );
  MUX2_X1 U448 ( .A(n219), .B(sll_14_ML_int_4__43_), .S(n206), .Z(
        sll_14_ML_int_5__59_) );
  MUX2_X1 U449 ( .A(n219), .B(n253), .S(n210), .Z(sll_14_ML_int_4__43_) );
  MUX2_X1 U450 ( .A(n218), .B(n259), .S(n213), .Z(n253) );
  MUX2_X1 U451 ( .A(n218), .B(sll_14_ML_int_4__44_), .S(n206), .Z(
        sll_14_ML_int_5__60_) );
  MUX2_X1 U452 ( .A(n218), .B(n254), .S(n210), .Z(sll_14_ML_int_4__44_) );
  MUX2_X1 U453 ( .A(n218), .B(n257), .S(n213), .Z(n254) );
  MUX2_X1 U454 ( .A(n218), .B(sll_14_ML_int_1__30_), .S(n216), .Z(n257) );
  MUX2_X1 U455 ( .A(n218), .B(sll_14_ML_int_4__45_), .S(n206), .Z(
        sll_14_ML_int_5__61_) );
  MUX2_X1 U456 ( .A(n218), .B(n255), .S(n210), .Z(sll_14_ML_int_4__45_) );
  MUX2_X1 U457 ( .A(n218), .B(n258), .S(n213), .Z(n255) );
  MUX2_X1 U458 ( .A(n218), .B(n260), .S(n215), .Z(n258) );
  MUX2_X1 U459 ( .A(n218), .B(sll_14_ML_int_5__31_), .S(n199), .Z(N69) );
  MUX2_X1 U460 ( .A(n249), .B(sll_14_ML_int_4__15_), .S(n204), .Z(
        sll_14_ML_int_5__31_) );
  MUX2_X1 U461 ( .A(n256), .B(sll_14_ML_int_3__23_), .S(n210), .Z(n249) );
  MUX2_X1 U462 ( .A(n259), .B(sll_14_ML_int_2__27_), .S(n213), .Z(n256) );
  MUX2_X1 U463 ( .A(n260), .B(sll_14_ML_int_1__29_), .S(n215), .Z(n259) );
  MUX2_X1 U464 ( .A(n218), .B(a[30]), .S(n66), .Z(n260) );
  XOR2_X1 U465 ( .A(add_30_carry[5]), .B(n199), .Z(N80) );
endmodule


module register_N64_1 ( clk, reset, reg_in, reg_out );
  input [63:0] reg_in;
  output [63:0] reg_out;
  input clk, reset;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73;

  SDFF_X1 reg_out_reg_63_ ( .D(1'b0), .SI(n65), .SE(reg_in[63]), .CK(clk), .Q(
        reg_out[63]) );
  SDFF_X1 reg_out_reg_62_ ( .D(1'b0), .SI(n65), .SE(reg_in[62]), .CK(clk), .Q(
        reg_out[62]) );
  SDFF_X1 reg_out_reg_61_ ( .D(1'b0), .SI(n65), .SE(reg_in[61]), .CK(clk), .Q(
        reg_out[61]) );
  SDFF_X1 reg_out_reg_60_ ( .D(1'b0), .SI(n65), .SE(reg_in[60]), .CK(clk), .Q(
        reg_out[60]) );
  SDFF_X1 reg_out_reg_59_ ( .D(1'b0), .SI(n65), .SE(reg_in[59]), .CK(clk), .Q(
        reg_out[59]) );
  SDFF_X1 reg_out_reg_58_ ( .D(1'b0), .SI(n65), .SE(reg_in[58]), .CK(clk), .Q(
        reg_out[58]) );
  SDFF_X1 reg_out_reg_57_ ( .D(1'b0), .SI(n65), .SE(reg_in[57]), .CK(clk), .Q(
        reg_out[57]) );
  SDFF_X1 reg_out_reg_56_ ( .D(1'b0), .SI(n65), .SE(reg_in[56]), .CK(clk), .Q(
        reg_out[56]) );
  SDFF_X1 reg_out_reg_55_ ( .D(1'b0), .SI(n65), .SE(reg_in[55]), .CK(clk), .Q(
        reg_out[55]) );
  SDFF_X1 reg_out_reg_54_ ( .D(1'b0), .SI(n65), .SE(reg_in[54]), .CK(clk), .Q(
        reg_out[54]) );
  SDFF_X1 reg_out_reg_53_ ( .D(1'b0), .SI(n65), .SE(reg_in[53]), .CK(clk), .Q(
        reg_out[53]) );
  SDFF_X1 reg_out_reg_52_ ( .D(1'b0), .SI(n66), .SE(reg_in[52]), .CK(clk), .Q(
        reg_out[52]) );
  SDFF_X1 reg_out_reg_51_ ( .D(1'b0), .SI(n66), .SE(reg_in[51]), .CK(clk), .Q(
        reg_out[51]) );
  SDFF_X1 reg_out_reg_50_ ( .D(1'b0), .SI(n66), .SE(reg_in[50]), .CK(clk), .Q(
        reg_out[50]) );
  SDFF_X1 reg_out_reg_49_ ( .D(1'b0), .SI(n66), .SE(reg_in[49]), .CK(clk), .Q(
        reg_out[49]) );
  SDFF_X1 reg_out_reg_48_ ( .D(1'b0), .SI(n66), .SE(reg_in[48]), .CK(clk), .Q(
        reg_out[48]) );
  SDFF_X1 reg_out_reg_47_ ( .D(1'b0), .SI(n66), .SE(reg_in[47]), .CK(clk), .Q(
        reg_out[47]) );
  SDFF_X1 reg_out_reg_46_ ( .D(1'b0), .SI(n66), .SE(reg_in[46]), .CK(clk), .Q(
        reg_out[46]) );
  SDFF_X1 reg_out_reg_45_ ( .D(1'b0), .SI(n66), .SE(reg_in[45]), .CK(clk), .Q(
        reg_out[45]) );
  SDFF_X1 reg_out_reg_44_ ( .D(1'b0), .SI(n66), .SE(reg_in[44]), .CK(clk), .Q(
        reg_out[44]) );
  SDFF_X1 reg_out_reg_43_ ( .D(1'b0), .SI(n66), .SE(reg_in[43]), .CK(clk), .Q(
        reg_out[43]) );
  SDFF_X1 reg_out_reg_42_ ( .D(1'b0), .SI(n66), .SE(reg_in[42]), .CK(clk), .Q(
        reg_out[42]) );
  SDFF_X1 reg_out_reg_41_ ( .D(1'b0), .SI(n67), .SE(reg_in[41]), .CK(clk), .Q(
        reg_out[41]) );
  SDFF_X1 reg_out_reg_40_ ( .D(1'b0), .SI(n67), .SE(reg_in[40]), .CK(clk), .Q(
        reg_out[40]) );
  SDFF_X1 reg_out_reg_39_ ( .D(1'b0), .SI(n67), .SE(reg_in[39]), .CK(clk), .Q(
        reg_out[39]) );
  SDFF_X1 reg_out_reg_38_ ( .D(1'b0), .SI(n67), .SE(reg_in[38]), .CK(clk), .Q(
        reg_out[38]) );
  SDFF_X1 reg_out_reg_37_ ( .D(1'b0), .SI(n67), .SE(reg_in[37]), .CK(clk), .Q(
        reg_out[37]) );
  SDFF_X1 reg_out_reg_36_ ( .D(1'b0), .SI(n67), .SE(reg_in[36]), .CK(clk), .Q(
        reg_out[36]) );
  SDFF_X1 reg_out_reg_35_ ( .D(1'b0), .SI(n67), .SE(reg_in[35]), .CK(clk), .Q(
        reg_out[35]) );
  SDFF_X1 reg_out_reg_34_ ( .D(1'b0), .SI(n67), .SE(reg_in[34]), .CK(clk), .Q(
        reg_out[34]) );
  SDFF_X1 reg_out_reg_33_ ( .D(1'b0), .SI(n67), .SE(reg_in[33]), .CK(clk), .Q(
        reg_out[33]) );
  SDFF_X1 reg_out_reg_32_ ( .D(1'b0), .SI(n67), .SE(reg_in[32]), .CK(clk), .Q(
        reg_out[32]) );
  SDFF_X1 reg_out_reg_31_ ( .D(1'b0), .SI(n67), .SE(reg_in[31]), .CK(clk), .Q(
        reg_out[31]) );
  SDFF_X1 reg_out_reg_30_ ( .D(1'b0), .SI(n68), .SE(reg_in[30]), .CK(clk), .Q(
        reg_out[30]) );
  SDFF_X1 reg_out_reg_29_ ( .D(1'b0), .SI(n68), .SE(reg_in[29]), .CK(clk), .Q(
        reg_out[29]) );
  SDFF_X1 reg_out_reg_28_ ( .D(1'b0), .SI(n68), .SE(reg_in[28]), .CK(clk), .Q(
        reg_out[28]) );
  SDFF_X1 reg_out_reg_27_ ( .D(1'b0), .SI(n68), .SE(reg_in[27]), .CK(clk), .Q(
        reg_out[27]) );
  SDFF_X1 reg_out_reg_26_ ( .D(1'b0), .SI(n68), .SE(reg_in[26]), .CK(clk), .Q(
        reg_out[26]) );
  SDFF_X1 reg_out_reg_25_ ( .D(1'b0), .SI(n68), .SE(reg_in[25]), .CK(clk), .Q(
        reg_out[25]) );
  SDFF_X1 reg_out_reg_24_ ( .D(1'b0), .SI(n68), .SE(reg_in[24]), .CK(clk), .Q(
        reg_out[24]) );
  SDFF_X1 reg_out_reg_23_ ( .D(1'b0), .SI(n68), .SE(reg_in[23]), .CK(clk), .Q(
        reg_out[23]) );
  SDFF_X1 reg_out_reg_22_ ( .D(1'b0), .SI(n68), .SE(reg_in[22]), .CK(clk), .Q(
        reg_out[22]) );
  SDFF_X1 reg_out_reg_21_ ( .D(1'b0), .SI(n68), .SE(reg_in[21]), .CK(clk), .Q(
        reg_out[21]) );
  SDFF_X1 reg_out_reg_20_ ( .D(1'b0), .SI(n68), .SE(reg_in[20]), .CK(clk), .Q(
        reg_out[20]) );
  SDFF_X1 reg_out_reg_19_ ( .D(1'b0), .SI(n69), .SE(reg_in[19]), .CK(clk), .Q(
        reg_out[19]) );
  SDFF_X1 reg_out_reg_18_ ( .D(1'b0), .SI(n69), .SE(reg_in[18]), .CK(clk), .Q(
        reg_out[18]) );
  SDFF_X1 reg_out_reg_17_ ( .D(1'b0), .SI(n69), .SE(reg_in[17]), .CK(clk), .Q(
        reg_out[17]) );
  SDFF_X1 reg_out_reg_16_ ( .D(1'b0), .SI(n69), .SE(reg_in[16]), .CK(clk), .Q(
        reg_out[16]) );
  SDFF_X1 reg_out_reg_15_ ( .D(1'b0), .SI(n69), .SE(reg_in[15]), .CK(clk), .Q(
        reg_out[15]) );
  SDFF_X1 reg_out_reg_14_ ( .D(1'b0), .SI(n69), .SE(reg_in[14]), .CK(clk), .Q(
        reg_out[14]) );
  SDFF_X1 reg_out_reg_13_ ( .D(1'b0), .SI(n69), .SE(reg_in[13]), .CK(clk), .Q(
        reg_out[13]) );
  SDFF_X1 reg_out_reg_12_ ( .D(1'b0), .SI(n69), .SE(reg_in[12]), .CK(clk), .Q(
        reg_out[12]) );
  SDFF_X1 reg_out_reg_11_ ( .D(1'b0), .SI(n69), .SE(reg_in[11]), .CK(clk), .Q(
        reg_out[11]) );
  SDFF_X1 reg_out_reg_10_ ( .D(1'b0), .SI(n69), .SE(reg_in[10]), .CK(clk), .Q(
        reg_out[10]) );
  SDFF_X1 reg_out_reg_9_ ( .D(1'b0), .SI(n69), .SE(reg_in[9]), .CK(clk), .Q(
        reg_out[9]) );
  SDFF_X1 reg_out_reg_8_ ( .D(1'b0), .SI(n70), .SE(reg_in[8]), .CK(clk), .Q(
        reg_out[8]) );
  SDFF_X1 reg_out_reg_7_ ( .D(1'b0), .SI(n70), .SE(reg_in[7]), .CK(clk), .Q(
        reg_out[7]) );
  SDFF_X1 reg_out_reg_6_ ( .D(1'b0), .SI(n70), .SE(reg_in[6]), .CK(clk), .Q(
        reg_out[6]) );
  SDFF_X1 reg_out_reg_5_ ( .D(1'b0), .SI(n70), .SE(reg_in[5]), .CK(clk), .Q(
        reg_out[5]) );
  SDFF_X1 reg_out_reg_4_ ( .D(1'b0), .SI(n70), .SE(reg_in[4]), .CK(clk), .Q(
        reg_out[4]) );
  SDFF_X1 reg_out_reg_3_ ( .D(1'b0), .SI(n70), .SE(reg_in[3]), .CK(clk), .Q(
        reg_out[3]) );
  SDFF_X1 reg_out_reg_2_ ( .D(1'b0), .SI(n70), .SE(reg_in[2]), .CK(clk), .Q(
        reg_out[2]) );
  SDFF_X1 reg_out_reg_1_ ( .D(1'b0), .SI(n70), .SE(reg_in[1]), .CK(clk), .Q(
        reg_out[1]) );
  SDFF_X1 reg_out_reg_0_ ( .D(1'b0), .SI(n70), .SE(reg_in[0]), .CK(clk), .Q(
        reg_out[0]) );
  BUF_X1 U67 ( .A(n71), .Z(n69) );
  BUF_X1 U68 ( .A(n71), .Z(n68) );
  BUF_X1 U69 ( .A(n72), .Z(n67) );
  BUF_X1 U70 ( .A(n72), .Z(n66) );
  BUF_X1 U71 ( .A(n72), .Z(n65) );
  BUF_X1 U72 ( .A(n71), .Z(n70) );
  INV_X1 U73 ( .A(reset), .ZN(n73) );
  BUF_X1 U74 ( .A(n73), .Z(n71) );
  BUF_X1 U75 ( .A(n73), .Z(n72) );
endmodule


module TopModule ( clk, iclk, a, b, reset, resetReg, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;
  input clk, iclk, reset, resetReg;

  wire   [31:0] mulA;
  wire   [31:0] mulB;
  wire   [63:0] mulResult;

  register_N64_0 R0 ( .clk(clk), .reset(resetReg), .reg_in({a, b}), .reg_out({
        mulA, mulB}) );
  sequentialMultiplier M0 ( .a(mulA), .b(mulB), .reset(reset), .clk(iclk), 
        .result(mulResult) );
  register_N64_1 R2 ( .clk(clk), .reset(resetReg), .reg_in(mulResult), 
        .reg_out(result) );
endmodule

