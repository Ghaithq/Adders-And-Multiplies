
module comparator8bit_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n4;
  wire   [7:4] carry;

  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(n1), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_3 ( .A(n4), .B(A[3]), .S(SUM[3]) );
  AND2_X1 U1 ( .A1(A[4]), .A2(carry[4]), .ZN(n1) );
  AND2_X1 U2 ( .A1(n4), .A2(A[3]), .ZN(carry[4]) );
  CLKBUF_X1 U3 ( .A(A[2]), .Z(n2) );
  XOR2_X1 U4 ( .A(A[1]), .B(A[0]), .Z(SUM[1]) );
  AND2_X1 U5 ( .A1(A[1]), .A2(A[0]), .ZN(n3) );
  AND2_X1 U6 ( .A1(A[2]), .A2(n3), .ZN(n4) );
  XOR2_X1 U7 ( .A(n2), .B(n3), .Z(SUM[2]) );
  XOR2_X1 U8 ( .A(carry[4]), .B(A[4]), .Z(SUM[4]) );
  XOR2_X1 U9 ( .A(carry[7]), .B(A[7]), .Z(SUM[7]) );
endmodule


module comparator8bit_DW01_add_2 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n28, n29, n30, n31, n32, n36, n37, n39,
         n40, n41, n42, n43, n45, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n91;

  OAI21_X1 U60 ( .B1(n12), .B2(n10), .A(n11), .ZN(SUM[8]) );
  OR2_X1 U61 ( .A1(B[0]), .A2(A[0]), .ZN(n81) );
  INV_X1 U62 ( .A(n86), .ZN(n28) );
  CLKBUF_X1 U63 ( .A(n21), .Z(n82) );
  BUF_X1 U64 ( .A(n32), .Z(n85) );
  CLKBUF_X1 U65 ( .A(n19), .Z(n83) );
  XNOR2_X1 U66 ( .A(n84), .B(n37), .ZN(SUM[1]) );
  NAND2_X1 U67 ( .A1(n36), .A2(n87), .ZN(n84) );
  AND2_X1 U68 ( .A1(B[3]), .A2(A[3]), .ZN(n86) );
  INV_X1 U69 ( .A(n88), .ZN(n36) );
  AND2_X1 U70 ( .A1(B[1]), .A2(A[1]), .ZN(n88) );
  OR2_X1 U71 ( .A1(B[1]), .A2(A[1]), .ZN(n87) );
  OAI21_X1 U72 ( .B1(n30), .B2(n85), .A(n31), .ZN(n89) );
  AND2_X1 U73 ( .A1(n81), .A2(n39), .ZN(SUM[0]) );
  INV_X1 U74 ( .A(n82), .ZN(n20) );
  XOR2_X1 U75 ( .A(n6), .B(n85), .Z(SUM[2]) );
  NAND2_X1 U76 ( .A1(n45), .A2(n31), .ZN(n6) );
  INV_X1 U77 ( .A(n30), .ZN(n45) );
  XOR2_X1 U78 ( .A(n24), .B(n4), .Z(SUM[4]) );
  NAND2_X1 U79 ( .A1(n43), .A2(n23), .ZN(n4) );
  INV_X1 U80 ( .A(n22), .ZN(n43) );
  OAI21_X1 U81 ( .B1(n32), .B2(n30), .A(n31), .ZN(n29) );
  INV_X1 U82 ( .A(n39), .ZN(n37) );
  XNOR2_X1 U83 ( .A(n5), .B(n89), .ZN(SUM[3]) );
  NAND2_X1 U84 ( .A1(n91), .A2(n28), .ZN(n5) );
  AOI21_X1 U85 ( .B1(n87), .B2(n37), .A(n88), .ZN(n32) );
  NAND2_X1 U86 ( .A1(n40), .A2(n11), .ZN(n1) );
  INV_X1 U87 ( .A(n10), .ZN(n40) );
  XOR2_X1 U88 ( .A(n3), .B(n20), .Z(SUM[5]) );
  NAND2_X1 U89 ( .A1(n42), .A2(n83), .ZN(n3) );
  INV_X1 U90 ( .A(n18), .ZN(n42) );
  XNOR2_X1 U91 ( .A(n2), .B(n17), .ZN(SUM[6]) );
  OAI21_X1 U92 ( .B1(n20), .B2(n18), .A(n83), .ZN(n17) );
  NAND2_X1 U93 ( .A1(B[2]), .A2(A[2]), .ZN(n31) );
  NOR2_X1 U94 ( .A1(A[5]), .A2(B[5]), .ZN(n18) );
  NOR2_X1 U95 ( .A1(B[2]), .A2(A[2]), .ZN(n30) );
  NOR2_X1 U96 ( .A1(B[6]), .A2(A[6]), .ZN(n15) );
  NAND2_X1 U97 ( .A1(B[4]), .A2(A[4]), .ZN(n23) );
  NOR2_X1 U98 ( .A1(B[4]), .A2(A[4]), .ZN(n22) );
  NAND2_X1 U99 ( .A1(B[7]), .A2(A[7]), .ZN(n11) );
  OR2_X1 U100 ( .A1(B[3]), .A2(A[3]), .ZN(n91) );
  NAND2_X1 U101 ( .A1(n41), .A2(n16), .ZN(n2) );
  INV_X1 U102 ( .A(n15), .ZN(n41) );
  NOR2_X1 U103 ( .A1(B[7]), .A2(A[7]), .ZN(n10) );
  NAND2_X1 U104 ( .A1(B[6]), .A2(A[6]), .ZN(n16) );
  NAND2_X1 U105 ( .A1(B[5]), .A2(A[5]), .ZN(n19) );
  OAI21_X1 U106 ( .B1(n24), .B2(n22), .A(n23), .ZN(n21) );
  AOI21_X1 U107 ( .B1(n29), .B2(n91), .A(n86), .ZN(n24) );
  NOR2_X1 U108 ( .A1(n15), .A2(n18), .ZN(n13) );
  AOI21_X1 U109 ( .B1(n13), .B2(n21), .A(n14), .ZN(n12) );
  XOR2_X1 U110 ( .A(n12), .B(n1), .Z(SUM[7]) );
  NAND2_X1 U111 ( .A1(B[0]), .A2(A[0]), .ZN(n39) );
  OAI21_X1 U112 ( .B1(n15), .B2(n19), .A(n16), .ZN(n14) );
endmodule


module comparator8bit ( a, b, f_bigger, diff );
  input [7:0] a;
  input [7:0] b;
  output [7:0] diff;
  output f_bigger;
  wire   temp_7_, temp_6_, temp_5_, temp_4_, temp_3_, temp_2_, temp_1_, N11,
         N12, N13, N14, N15, N16, N17, complement_b_7_, complement_b_6_,
         complement_b_5_, complement_b_4_, complement_b_3_, complement_b_2_,
         complement_b_1_, n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         SYNOPSYS_UNCONNECTED_1;

  comparator8bit_DW01_inc_0 add_18 ( .A({n21, n22, n23, n24, n25, n26, n27, 
        n18}), .SUM({N17, N16, N15, N14, N13, N12, N11, SYNOPSYS_UNCONNECTED_1}) );
  comparator8bit_DW01_add_2 add_14 ( .A({1'b0, a}), .B({1'b0, complement_b_7_, 
        complement_b_6_, complement_b_5_, complement_b_4_, complement_b_3_, 
        complement_b_2_, complement_b_1_, n2}), .CI(1'b0), .SUM({f_bigger, 
        temp_7_, temp_6_, temp_5_, temp_4_, temp_3_, temp_2_, temp_1_, diff[0]}) );
  MUX2_X1 U3 ( .A(N11), .B(temp_1_), .S(n9), .Z(diff[1]) );
  NOR3_X1 U5 ( .A1(n7), .A2(n16), .A3(n14), .ZN(n11) );
  OR3_X1 U6 ( .A1(b[1]), .A2(b[2]), .A3(b[4]), .ZN(n13) );
  BUF_X1 U7 ( .A(b[0]), .Z(n2) );
  OR2_X1 U8 ( .A1(b[1]), .A2(b[2]), .ZN(n1) );
  MUX2_X1 U9 ( .A(temp_3_), .B(N13), .S(n8), .Z(diff[3]) );
  XNOR2_X1 U10 ( .A(n3), .B(b[3]), .ZN(complement_b_3_) );
  NOR2_X1 U11 ( .A1(n1), .A2(n2), .ZN(n3) );
  MUX2_X2 U12 ( .A(N12), .B(temp_2_), .S(n9), .Z(diff[2]) );
  XNOR2_X1 U13 ( .A(n4), .B(b[5]), .ZN(complement_b_5_) );
  NOR2_X1 U14 ( .A1(n13), .A2(n14), .ZN(n4) );
  CLKBUF_X1 U15 ( .A(b[2]), .Z(n5) );
  OR2_X1 U16 ( .A1(b[1]), .A2(b[2]), .ZN(n7) );
  MUX2_X1 U17 ( .A(N14), .B(temp_4_), .S(n17), .Z(diff[4]) );
  INV_X1 U18 ( .A(n17), .ZN(n8) );
  INV_X1 U19 ( .A(n8), .ZN(n9) );
  OR2_X1 U20 ( .A1(n13), .A2(n14), .ZN(n10) );
  XNOR2_X1 U21 ( .A(n11), .B(b[6]), .ZN(complement_b_6_) );
  CLKBUF_X1 U22 ( .A(f_bigger), .Z(n17) );
  OR2_X1 U23 ( .A1(n14), .A2(n7), .ZN(n19) );
  OR2_X1 U24 ( .A1(b[6]), .A2(b[5]), .ZN(n12) );
  OR2_X1 U25 ( .A1(b[0]), .A2(b[3]), .ZN(n14) );
  XNOR2_X1 U26 ( .A(n15), .B(b[7]), .ZN(complement_b_7_) );
  NOR2_X1 U27 ( .A1(n10), .A2(n12), .ZN(n15) );
  OR2_X1 U28 ( .A1(b[5]), .A2(b[4]), .ZN(n16) );
  OR2_X1 U29 ( .A1(b[1]), .A2(b[0]), .ZN(n20) );
  INV_X1 U30 ( .A(diff[0]), .ZN(n18) );
  XOR2_X1 U31 ( .A(n19), .B(b[4]), .Z(complement_b_4_) );
  XOR2_X1 U32 ( .A(n20), .B(n5), .Z(complement_b_2_) );
  XOR2_X1 U33 ( .A(b[1]), .B(b[0]), .Z(complement_b_1_) );
  INV_X1 U34 ( .A(temp_7_), .ZN(n21) );
  INV_X1 U35 ( .A(temp_6_), .ZN(n22) );
  INV_X1 U36 ( .A(temp_5_), .ZN(n23) );
  INV_X1 U37 ( .A(temp_4_), .ZN(n24) );
  INV_X1 U38 ( .A(temp_3_), .ZN(n25) );
  INV_X1 U39 ( .A(temp_2_), .ZN(n26) );
  INV_X1 U40 ( .A(temp_1_), .ZN(n27) );
  MUX2_X1 U41 ( .A(N15), .B(temp_5_), .S(n9), .Z(diff[5]) );
  MUX2_X1 U42 ( .A(N16), .B(temp_6_), .S(n9), .Z(diff[6]) );
  MUX2_X1 U43 ( .A(N17), .B(temp_7_), .S(n9), .Z(diff[7]) );
endmodule


module shiftRegister_DW_rightsh_2 ( A, DATA_TC, SH, B );
  input [23:0] A;
  input [4:0] SH;
  output [23:0] B;
  input DATA_TC;
  wire   n1, n3, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248;

  INV_X1 U155 ( .A(n248), .ZN(n246) );
  MUX2_X1 U156 ( .A(n12), .B(n14), .S(SH[1]), .Z(B[5]) );
  MUX2_X1 U157 ( .A(n8), .B(n10), .S(SH[1]), .Z(B[1]) );
  MUX2_X1 U158 ( .A(n9), .B(n7), .S(n1), .Z(B[0]) );
  MUX2_X1 U159 ( .A(n25), .B(n27), .S(SH[1]), .Z(B[18]) );
  MUX2_X1 U160 ( .A(n28), .B(n30), .S(SH[1]), .Z(B[21]) );
  MUX2_X1 U161 ( .A(n27), .B(n29), .S(SH[1]), .Z(B[20]) );
  BUF_X1 U162 ( .A(SH[3]), .Z(n197) );
  INV_X1 U163 ( .A(n248), .ZN(n247) );
  NAND2_X1 U164 ( .A1(A[17]), .A2(SH[0]), .ZN(n225) );
  NAND2_X1 U165 ( .A1(A[2]), .A2(n208), .ZN(n187) );
  NAND2_X1 U166 ( .A1(A[3]), .A2(n247), .ZN(n188) );
  NAND2_X1 U167 ( .A1(n187), .A2(n188), .ZN(n106) );
  INV_X2 U168 ( .A(n244), .ZN(n63) );
  NAND2_X1 U169 ( .A1(n49), .A2(n3), .ZN(n189) );
  NAND2_X1 U170 ( .A1(n53), .A2(SH[2]), .ZN(n190) );
  NAND2_X1 U171 ( .A1(n189), .A2(n190), .ZN(n17) );
  BUF_X1 U172 ( .A(SH[4]), .Z(n244) );
  NAND2_X1 U173 ( .A1(A[19]), .A2(n191), .ZN(n192) );
  NAND2_X1 U174 ( .A1(A[20]), .A2(n246), .ZN(n193) );
  NAND2_X1 U175 ( .A1(n192), .A2(n193), .ZN(n123) );
  INV_X1 U176 ( .A(n246), .ZN(n191) );
  NAND2_X1 U177 ( .A1(n109), .A2(n194), .ZN(n195) );
  NAND2_X1 U178 ( .A1(n245), .A2(n125), .ZN(n196) );
  NAND2_X1 U179 ( .A1(n195), .A2(n196), .ZN(n84) );
  INV_X1 U180 ( .A(n245), .ZN(n194) );
  BUF_X2 U181 ( .A(SH[4]), .Z(n245) );
  BUF_X2 U182 ( .A(SH[3]), .Z(n199) );
  BUF_X2 U183 ( .A(SH[3]), .Z(n198) );
  NAND2_X1 U184 ( .A1(A[1]), .A2(n200), .ZN(n201) );
  NAND2_X1 U185 ( .A1(A[0]), .A2(n248), .ZN(n202) );
  NAND2_X1 U186 ( .A1(n201), .A2(n202), .ZN(n104) );
  INV_X1 U187 ( .A(n248), .ZN(n200) );
  NAND2_X1 U188 ( .A1(A[7]), .A2(n200), .ZN(n203) );
  NAND2_X1 U189 ( .A1(A[6]), .A2(n248), .ZN(n204) );
  NAND2_X1 U190 ( .A1(n204), .A2(n203), .ZN(n110) );
  NAND2_X1 U191 ( .A1(A[20]), .A2(n205), .ZN(n206) );
  NAND2_X1 U192 ( .A1(A[21]), .A2(n246), .ZN(n207) );
  NAND2_X1 U193 ( .A1(n206), .A2(n207), .ZN(n124) );
  INV_X1 U194 ( .A(n246), .ZN(n205) );
  NAND2_X1 U195 ( .A1(A[18]), .A2(n208), .ZN(n209) );
  NAND2_X1 U196 ( .A1(A[19]), .A2(n246), .ZN(n210) );
  NAND2_X1 U197 ( .A1(n209), .A2(n210), .ZN(n122) );
  INV_X1 U198 ( .A(n246), .ZN(n208) );
  NAND2_X1 U199 ( .A1(A[17]), .A2(n211), .ZN(n212) );
  NAND2_X1 U200 ( .A1(A[18]), .A2(n246), .ZN(n213) );
  NAND2_X1 U201 ( .A1(n212), .A2(n213), .ZN(n121) );
  INV_X1 U202 ( .A(n246), .ZN(n211) );
  NAND2_X1 U203 ( .A1(n82), .A2(n214), .ZN(n215) );
  NAND2_X1 U204 ( .A1(n90), .A2(n199), .ZN(n216) );
  NAND2_X1 U205 ( .A1(n215), .A2(n216), .ZN(n42) );
  INV_X1 U206 ( .A(n198), .ZN(n214) );
  NAND2_X1 U207 ( .A1(n86), .A2(n228), .ZN(n217) );
  NAND2_X1 U208 ( .A1(n94), .A2(n199), .ZN(n218) );
  NAND2_X1 U209 ( .A1(n217), .A2(n218), .ZN(n46) );
  NAND2_X1 U210 ( .A1(n84), .A2(n219), .ZN(n220) );
  NAND2_X1 U211 ( .A1(n92), .A2(n198), .ZN(n221) );
  NAND2_X1 U212 ( .A1(n220), .A2(n221), .ZN(n44) );
  INV_X1 U213 ( .A(n198), .ZN(n219) );
  NAND2_X1 U214 ( .A1(n93), .A2(n219), .ZN(n222) );
  NAND2_X1 U215 ( .A1(n101), .A2(n198), .ZN(n223) );
  NAND2_X1 U216 ( .A1(n223), .A2(n222), .ZN(n53) );
  MUX2_X1 U217 ( .A(A[22]), .B(A[21]), .S(n248), .Z(n125) );
  NAND2_X1 U218 ( .A1(A[16]), .A2(n191), .ZN(n224) );
  NAND2_X1 U219 ( .A1(n225), .A2(n224), .ZN(n120) );
  NAND2_X1 U220 ( .A1(A[22]), .A2(n205), .ZN(n226) );
  NAND2_X1 U221 ( .A1(A[23]), .A2(n246), .ZN(n227) );
  NAND2_X1 U222 ( .A1(n226), .A2(n227), .ZN(n126) );
  NAND2_X1 U223 ( .A1(n83), .A2(n228), .ZN(n229) );
  NAND2_X1 U224 ( .A1(n91), .A2(n199), .ZN(n230) );
  NAND2_X1 U225 ( .A1(n229), .A2(n230), .ZN(n43) );
  INV_X1 U226 ( .A(n197), .ZN(n228) );
  NAND2_X1 U227 ( .A1(n194), .A2(n106), .ZN(n231) );
  NAND2_X1 U228 ( .A1(n122), .A2(n245), .ZN(n232) );
  NAND2_X1 U229 ( .A1(n232), .A2(n231), .ZN(n81) );
  NAND2_X1 U230 ( .A1(n104), .A2(n63), .ZN(n233) );
  NAND2_X1 U231 ( .A1(n120), .A2(n245), .ZN(n234) );
  NAND2_X1 U232 ( .A1(n234), .A2(n233), .ZN(n79) );
  NAND2_X1 U233 ( .A1(n110), .A2(n63), .ZN(n236) );
  NAND2_X1 U234 ( .A1(n126), .A2(n245), .ZN(n237) );
  NAND2_X1 U235 ( .A1(n237), .A2(n236), .ZN(n85) );
  INV_X1 U236 ( .A(n245), .ZN(n235) );
  NAND2_X1 U237 ( .A1(n108), .A2(n235), .ZN(n238) );
  NAND2_X1 U238 ( .A1(n124), .A2(n245), .ZN(n239) );
  NAND2_X1 U239 ( .A1(n238), .A2(n239), .ZN(n83) );
  NAND2_X1 U240 ( .A1(n81), .A2(n228), .ZN(n240) );
  NAND2_X1 U241 ( .A1(n89), .A2(n198), .ZN(n241) );
  NAND2_X1 U242 ( .A1(n240), .A2(n241), .ZN(n41) );
  NAND2_X1 U243 ( .A1(n85), .A2(n228), .ZN(n242) );
  NAND2_X1 U244 ( .A1(n93), .A2(n198), .ZN(n243) );
  NAND2_X1 U245 ( .A1(n242), .A2(n243), .ZN(n45) );
  AND2_X1 U246 ( .A1(n29), .A2(n1), .ZN(B[22]) );
  AND2_X1 U247 ( .A1(n30), .A2(n1), .ZN(B[23]) );
  AND2_X1 U248 ( .A1(n61), .A2(n3), .ZN(n29) );
  AND2_X1 U249 ( .A1(n62), .A2(n3), .ZN(n30) );
  AND2_X1 U250 ( .A1(n60), .A2(n3), .ZN(n28) );
  AND2_X1 U251 ( .A1(n59), .A2(n3), .ZN(n27) );
  INV_X1 U252 ( .A(n197), .ZN(n31) );
  INV_X1 U253 ( .A(SH[2]), .ZN(n3) );
  INV_X1 U254 ( .A(SH[1]), .ZN(n1) );
  MUX2_X1 U255 ( .A(n21), .B(n23), .S(SH[1]), .Z(B[14]) );
  MUX2_X1 U256 ( .A(n23), .B(n25), .S(SH[1]), .Z(B[16]) );
  MUX2_X1 U257 ( .A(n26), .B(n28), .S(SH[1]), .Z(B[19]) );
  MUX2_X1 U258 ( .A(n24), .B(n26), .S(SH[1]), .Z(B[17]) );
  MUX2_X1 U259 ( .A(n22), .B(n24), .S(SH[1]), .Z(B[15]) );
  MUX2_X1 U260 ( .A(n17), .B(n19), .S(SH[1]), .Z(B[10]) );
  MUX2_X1 U261 ( .A(n11), .B(n13), .S(SH[1]), .Z(B[4]) );
  MUX2_X1 U262 ( .A(n15), .B(n17), .S(SH[1]), .Z(B[8]) );
  MUX2_X1 U263 ( .A(n13), .B(n15), .S(SH[1]), .Z(B[6]) );
  MUX2_X1 U264 ( .A(n14), .B(n16), .S(SH[1]), .Z(B[7]) );
  MUX2_X1 U265 ( .A(n20), .B(n22), .S(SH[1]), .Z(B[13]) );
  MUX2_X1 U266 ( .A(n57), .B(n61), .S(SH[2]), .Z(n25) );
  MUX2_X1 U267 ( .A(n58), .B(n62), .S(SH[2]), .Z(n26) );
  MUX2_X1 U268 ( .A(n47), .B(n51), .S(SH[2]), .Z(n15) );
  MUX2_X1 U269 ( .A(n55), .B(n59), .S(SH[2]), .Z(n23) );
  MUX2_X1 U270 ( .A(n56), .B(n60), .S(SH[2]), .Z(n24) );
  MUX2_X1 U271 ( .A(n54), .B(n58), .S(SH[2]), .Z(n22) );
  MUX2_X1 U272 ( .A(n51), .B(n55), .S(SH[2]), .Z(n19) );
  MUX2_X1 U273 ( .A(n48), .B(n52), .S(SH[2]), .Z(n16) );
  MUX2_X1 U274 ( .A(n53), .B(n57), .S(SH[2]), .Z(n21) );
  MUX2_X1 U275 ( .A(n52), .B(n56), .S(SH[2]), .Z(n20) );
  MUX2_X1 U276 ( .A(n50), .B(n54), .S(SH[2]), .Z(n18) );
  AND2_X1 U277 ( .A1(n101), .A2(n31), .ZN(n61) );
  AND2_X1 U278 ( .A1(n102), .A2(n31), .ZN(n62) );
  AND2_X1 U279 ( .A1(n100), .A2(n31), .ZN(n60) );
  AND2_X1 U280 ( .A1(n99), .A2(n31), .ZN(n59) );
  AND2_X1 U281 ( .A1(n97), .A2(n31), .ZN(n57) );
  AND2_X1 U282 ( .A1(n98), .A2(n31), .ZN(n58) );
  AND2_X1 U283 ( .A1(n95), .A2(n31), .ZN(n55) );
  AND2_X1 U284 ( .A1(n96), .A2(n31), .ZN(n56) );
  MUX2_X1 U285 ( .A(n10), .B(n12), .S(SH[1]), .Z(B[3]) );
  MUX2_X1 U286 ( .A(n40), .B(n44), .S(SH[2]), .Z(n8) );
  MUX2_X1 U287 ( .A(n80), .B(n88), .S(n198), .Z(n40) );
  MUX2_X1 U288 ( .A(n105), .B(n121), .S(n245), .Z(n80) );
  MUX2_X1 U289 ( .A(n46), .B(n50), .S(SH[2]), .Z(n14) );
  MUX2_X1 U290 ( .A(n44), .B(n48), .S(SH[2]), .Z(n12) );
  MUX2_X1 U291 ( .A(n91), .B(n99), .S(n199), .Z(n51) );
  MUX2_X1 U292 ( .A(n92), .B(n100), .S(n199), .Z(n52) );
  MUX2_X1 U293 ( .A(n90), .B(n98), .S(n199), .Z(n50) );
  MUX2_X1 U294 ( .A(n88), .B(n96), .S(n198), .Z(n48) );
  MUX2_X1 U295 ( .A(n94), .B(n102), .S(n198), .Z(n54) );
  MUX2_X1 U296 ( .A(n89), .B(n97), .S(n198), .Z(n49) );
  MUX2_X1 U297 ( .A(n87), .B(n95), .S(n199), .Z(n47) );
  AND2_X1 U298 ( .A1(n127), .A2(n63), .ZN(n102) );
  AND2_X1 U299 ( .A1(n124), .A2(n63), .ZN(n99) );
  AND2_X1 U300 ( .A1(n122), .A2(n63), .ZN(n97) );
  AND2_X1 U301 ( .A1(n120), .A2(n63), .ZN(n95) );
  AND2_X1 U302 ( .A1(n123), .A2(n63), .ZN(n98) );
  AND2_X1 U303 ( .A1(n121), .A2(n63), .ZN(n96) );
  MUX2_X1 U304 ( .A(n39), .B(n43), .S(SH[2]), .Z(n7) );
  MUX2_X1 U305 ( .A(n79), .B(n87), .S(n198), .Z(n39) );
  MUX2_X1 U306 ( .A(A[5]), .B(A[6]), .S(n247), .Z(n109) );
  MUX2_X1 U307 ( .A(A[4]), .B(A[5]), .S(n247), .Z(n108) );
  MUX2_X1 U308 ( .A(A[14]), .B(A[15]), .S(n246), .Z(n118) );
  AND2_X1 U309 ( .A1(n112), .A2(n63), .ZN(n87) );
  MUX2_X1 U310 ( .A(A[8]), .B(A[9]), .S(n247), .Z(n112) );
  AND2_X1 U311 ( .A1(n116), .A2(n235), .ZN(n91) );
  MUX2_X1 U312 ( .A(A[12]), .B(A[13]), .S(n246), .Z(n116) );
  AND2_X1 U313 ( .A1(n113), .A2(n63), .ZN(n88) );
  MUX2_X1 U314 ( .A(A[9]), .B(A[10]), .S(n247), .Z(n113) );
  AND2_X1 U315 ( .A1(n117), .A2(n63), .ZN(n92) );
  MUX2_X1 U316 ( .A(A[13]), .B(A[14]), .S(n246), .Z(n117) );
  AND2_X1 U317 ( .A1(n115), .A2(n63), .ZN(n90) );
  MUX2_X1 U318 ( .A(A[11]), .B(A[12]), .S(n246), .Z(n115) );
  AND2_X1 U319 ( .A1(n119), .A2(n63), .ZN(n94) );
  MUX2_X1 U320 ( .A(A[15]), .B(A[16]), .S(n246), .Z(n119) );
  AND2_X1 U321 ( .A1(A[23]), .A2(n248), .ZN(n127) );
  MUX2_X1 U322 ( .A(n42), .B(n46), .S(SH[2]), .Z(n10) );
  MUX2_X1 U323 ( .A(n107), .B(n123), .S(n245), .Z(n82) );
  MUX2_X1 U324 ( .A(A[3]), .B(A[4]), .S(n247), .Z(n107) );
  MUX2_X1 U325 ( .A(n111), .B(n127), .S(n245), .Z(n86) );
  MUX2_X1 U326 ( .A(A[7]), .B(A[8]), .S(n247), .Z(n111) );
  MUX2_X1 U327 ( .A(A[1]), .B(A[2]), .S(n247), .Z(n105) );
  AND2_X1 U328 ( .A1(n114), .A2(n235), .ZN(n89) );
  MUX2_X1 U329 ( .A(A[10]), .B(A[11]), .S(n247), .Z(n114) );
  AND2_X1 U330 ( .A1(n118), .A2(n235), .ZN(n93) );
  MUX2_X1 U331 ( .A(n19), .B(n21), .S(SH[1]), .Z(B[12]) );
  AND2_X1 U332 ( .A1(n125), .A2(n63), .ZN(n100) );
  MUX2_X1 U333 ( .A(n18), .B(n20), .S(SH[1]), .Z(B[11]) );
  MUX2_X1 U334 ( .A(n16), .B(n18), .S(SH[1]), .Z(B[9]) );
  AND2_X1 U335 ( .A1(n126), .A2(n63), .ZN(n101) );
  MUX2_X1 U336 ( .A(n45), .B(n49), .S(SH[2]), .Z(n13) );
  MUX2_X1 U337 ( .A(n9), .B(n11), .S(SH[1]), .Z(B[2]) );
  MUX2_X1 U338 ( .A(n41), .B(n45), .S(SH[2]), .Z(n9) );
  MUX2_X1 U339 ( .A(n43), .B(n47), .S(SH[2]), .Z(n11) );
  INV_X1 U340 ( .A(SH[0]), .ZN(n248) );
endmodule


module shiftRegister ( a, b, f_bigger, shiftAmount, shiftedResult );
  input [23:0] a;
  input [23:0] b;
  input [4:0] shiftAmount;
  output [23:0] shiftedResult;
  input f_bigger;
  wire   n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  shiftRegister_DW_rightsh_2 srl_15 ( .A({n11, n12, n13, n14, n16, n17, n18, 
        n19, n20, n21, n22, n23, n24, n25, n2, n4, n5, n6, n7, n8, n9, n10, 
        n15, n26}), .DATA_TC(1'b0), .SH(shiftAmount), .B(shiftedResult) );
  CLKBUF_X1 U2 ( .A(f_bigger), .Z(n1) );
  MUX2_X1 U3 ( .A(a[23]), .B(b[23]), .S(n1), .Z(n11) );
  MUX2_X1 U4 ( .A(a[22]), .B(b[22]), .S(f_bigger), .Z(n12) );
  MUX2_X1 U5 ( .A(a[21]), .B(b[21]), .S(f_bigger), .Z(n13) );
  MUX2_X1 U6 ( .A(a[20]), .B(b[20]), .S(f_bigger), .Z(n14) );
  MUX2_X1 U7 ( .A(a[19]), .B(b[19]), .S(f_bigger), .Z(n16) );
  MUX2_X1 U8 ( .A(a[18]), .B(b[18]), .S(f_bigger), .Z(n17) );
  MUX2_X1 U9 ( .A(a[17]), .B(b[17]), .S(f_bigger), .Z(n18) );
  MUX2_X1 U10 ( .A(a[16]), .B(b[16]), .S(f_bigger), .Z(n19) );
  MUX2_X1 U11 ( .A(a[15]), .B(b[15]), .S(f_bigger), .Z(n20) );
  MUX2_X1 U12 ( .A(a[14]), .B(b[14]), .S(f_bigger), .Z(n21) );
  MUX2_X1 U13 ( .A(a[13]), .B(b[13]), .S(f_bigger), .Z(n22) );
  MUX2_X1 U14 ( .A(a[12]), .B(b[12]), .S(f_bigger), .Z(n23) );
  MUX2_X1 U15 ( .A(a[11]), .B(b[11]), .S(f_bigger), .Z(n24) );
  MUX2_X1 U16 ( .A(a[10]), .B(b[10]), .S(f_bigger), .Z(n25) );
  MUX2_X1 U17 ( .A(a[9]), .B(b[9]), .S(f_bigger), .Z(n2) );
  MUX2_X1 U18 ( .A(a[8]), .B(b[8]), .S(f_bigger), .Z(n4) );
  MUX2_X1 U19 ( .A(a[7]), .B(b[7]), .S(f_bigger), .Z(n5) );
  MUX2_X1 U20 ( .A(a[6]), .B(b[6]), .S(f_bigger), .Z(n6) );
  MUX2_X1 U21 ( .A(a[5]), .B(b[5]), .S(f_bigger), .Z(n7) );
  MUX2_X1 U22 ( .A(a[4]), .B(b[4]), .S(f_bigger), .Z(n8) );
  MUX2_X1 U23 ( .A(a[3]), .B(b[3]), .S(f_bigger), .Z(n9) );
  MUX2_X1 U24 ( .A(a[2]), .B(b[2]), .S(f_bigger), .Z(n10) );
  MUX2_X1 U25 ( .A(a[1]), .B(b[1]), .S(f_bigger), .Z(n15) );
  MUX2_X1 U26 ( .A(a[0]), .B(b[0]), .S(f_bigger), .Z(n26) );
endmodule


module carryLookAheadAdder ( a, b, cin, result, cout );
  input [23:0] a;
  input [23:0] b;
  output [23:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153;

  INV_X1 U1 ( .A(n1), .ZN(n144) );
  XOR2_X1 U2 ( .A(a[18]), .B(b[18]), .Z(n1) );
  NAND2_X1 U3 ( .A1(n100), .A2(n3), .ZN(n4) );
  NAND2_X1 U4 ( .A1(n2), .A2(b[20]), .ZN(n5) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(n147) );
  INV_X1 U6 ( .A(n100), .ZN(n2) );
  INV_X1 U7 ( .A(b[20]), .ZN(n3) );
  OAI22_X1 U8 ( .A1(n149), .A2(n17), .B1(n102), .B2(n101), .ZN(n28) );
  AOI22_X1 U9 ( .A1(a[21]), .A2(b[21]), .B1(n150), .B2(n6), .ZN(n103) );
  INV_X1 U10 ( .A(n149), .ZN(n6) );
  XNOR2_X1 U11 ( .A(a[13]), .B(b[13]), .ZN(n136) );
  AOI22_X1 U12 ( .A1(a[15]), .A2(b[15]), .B1(n13), .B2(n140), .ZN(n14) );
  XNOR2_X1 U13 ( .A(a[15]), .B(b[15]), .ZN(n139) );
  OAI22_X1 U14 ( .A1(n10), .A2(n135), .B1(n83), .B2(n82), .ZN(n137) );
  XNOR2_X1 U15 ( .A(a[9]), .B(b[9]), .ZN(n130) );
  OAI22_X1 U16 ( .A1(n12), .A2(n138), .B1(n87), .B2(n86), .ZN(n140) );
  AOI22_X1 U17 ( .A1(a[9]), .A2(b[9]), .B1(n131), .B2(n7), .ZN(n8) );
  INV_X1 U18 ( .A(n130), .ZN(n7) );
  AOI22_X1 U19 ( .A1(a[11]), .A2(b[11]), .B1(n134), .B2(n9), .ZN(n10) );
  INV_X1 U20 ( .A(n133), .ZN(n9) );
  AOI22_X1 U21 ( .A1(a[13]), .A2(b[13]), .B1(n137), .B2(n11), .ZN(n12) );
  INV_X1 U22 ( .A(n136), .ZN(n11) );
  INV_X1 U23 ( .A(n139), .ZN(n13) );
  AOI22_X1 U24 ( .A1(a[18]), .A2(b[18]), .B1(n145), .B2(n1), .ZN(n15) );
  AOI22_X1 U25 ( .A1(a[20]), .A2(b[20]), .B1(n148), .B2(n16), .ZN(n17) );
  INV_X1 U26 ( .A(n147), .ZN(n16) );
  INV_X1 U27 ( .A(n17), .ZN(n150) );
  INV_X1 U28 ( .A(n115), .ZN(n18) );
  INV_X1 U29 ( .A(n29), .ZN(n19) );
  INV_X1 U30 ( .A(n39), .ZN(n20) );
  INV_X1 U31 ( .A(n36), .ZN(n21) );
  CLKBUF_X1 U32 ( .A(n8), .Z(n22) );
  INV_X1 U33 ( .A(n41), .ZN(n23) );
  INV_X1 U34 ( .A(n32), .ZN(n24) );
  XNOR2_X1 U35 ( .A(a[2]), .B(b[2]), .ZN(n113) );
  INV_X1 U36 ( .A(n38), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n59), .A2(n58), .B1(n116), .B2(n24), .ZN(n26) );
  INV_X1 U38 ( .A(n45), .ZN(n27) );
  OAI22_X1 U39 ( .A1(n91), .A2(n90), .B1(n141), .B2(n14), .ZN(n29) );
  OAI22_X1 U40 ( .A1(n71), .A2(n70), .B1(n126), .B2(n20), .ZN(n30) );
  INV_X1 U41 ( .A(n18), .ZN(n31) );
  OAI22_X1 U42 ( .A1(n56), .A2(n55), .B1(n113), .B2(n18), .ZN(n32) );
  OAI22_X1 U43 ( .A1(n98), .A2(n97), .B1(n146), .B2(n15), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n100), .A2(n3), .B1(n147), .B2(n99), .ZN(n34) );
  OAI22_X1 U45 ( .A1(n85), .A2(n84), .B1(n136), .B2(n25), .ZN(n35) );
  OAI22_X1 U46 ( .A1(n87), .A2(n86), .B1(n138), .B2(n12), .ZN(n36) );
  OAI22_X1 U47 ( .A1(n78), .A2(n77), .B1(n132), .B2(n22), .ZN(n37) );
  OAI22_X1 U48 ( .A1(n83), .A2(n82), .B1(n135), .B2(n10), .ZN(n38) );
  OAI22_X1 U49 ( .A1(n68), .A2(n67), .B1(n124), .B2(n66), .ZN(n39) );
  OAI22_X1 U50 ( .A1(n105), .A2(n104), .B1(n103), .B2(n151), .ZN(n40) );
  OAI22_X1 U51 ( .A1(n94), .A2(n93), .B1(n142), .B2(n19), .ZN(n41) );
  OAI22_X1 U52 ( .A1(n81), .A2(n80), .B1(n133), .B2(n79), .ZN(n42) );
  OAI22_X1 U53 ( .A1(n62), .A2(n61), .B1(n119), .B2(n60), .ZN(n43) );
  OAI22_X1 U54 ( .A1(n65), .A2(n64), .B1(n122), .B2(n63), .ZN(n44) );
  OAI22_X1 U55 ( .A1(n74), .A2(n73), .B1(n128), .B2(n72), .ZN(n45) );
  OAI22_X1 U56 ( .A1(n89), .A2(n88), .B1(n139), .B2(n21), .ZN(n46) );
  XNOR2_X1 U57 ( .A(n34), .B(n149), .ZN(result[21]) );
  XNOR2_X1 U58 ( .A(n33), .B(n147), .ZN(result[20]) );
  XNOR2_X1 U59 ( .A(n47), .B(n146), .ZN(result[19]) );
  XNOR2_X1 U60 ( .A(n41), .B(n144), .ZN(result[18]) );
  XNOR2_X1 U61 ( .A(n29), .B(n142), .ZN(result[17]) );
  XNOR2_X1 U62 ( .A(n46), .B(n141), .ZN(result[16]) );
  XNOR2_X1 U63 ( .A(n36), .B(n139), .ZN(result[15]) );
  XNOR2_X1 U64 ( .A(n35), .B(n138), .ZN(result[14]) );
  XNOR2_X1 U65 ( .A(n38), .B(n136), .ZN(result[13]) );
  XNOR2_X1 U66 ( .A(n42), .B(n135), .ZN(result[12]) );
  XNOR2_X1 U67 ( .A(n37), .B(n133), .ZN(result[11]) );
  XNOR2_X1 U68 ( .A(n48), .B(n132), .ZN(result[10]) );
  XNOR2_X1 U69 ( .A(n45), .B(n130), .ZN(result[9]) );
  XNOR2_X1 U70 ( .A(n30), .B(n128), .ZN(result[8]) );
  XNOR2_X1 U71 ( .A(n43), .B(n122), .ZN(result[5]) );
  XNOR2_X1 U72 ( .A(n44), .B(n124), .ZN(result[6]) );
  XNOR2_X1 U73 ( .A(n39), .B(n126), .ZN(result[7]) );
  XNOR2_X1 U74 ( .A(n28), .B(n151), .ZN(result[22]) );
  XNOR2_X1 U75 ( .A(n153), .B(n152), .ZN(result[23]) );
  XNOR2_X1 U76 ( .A(cin), .B(n109), .ZN(result[0]) );
  OAI22_X1 U77 ( .A1(n96), .A2(n95), .B1(n144), .B2(n23), .ZN(n47) );
  OAI22_X1 U78 ( .A1(n76), .A2(n75), .B1(n130), .B2(n27), .ZN(n48) );
  XNOR2_X1 U79 ( .A(b[1]), .B(a[1]), .ZN(n110) );
  INV_X1 U80 ( .A(a[23]), .ZN(n107) );
  XOR2_X1 U81 ( .A(n107), .B(b[23]), .Z(n152) );
  INV_X1 U82 ( .A(a[22]), .ZN(n105) );
  INV_X1 U83 ( .A(b[22]), .ZN(n104) );
  XOR2_X1 U84 ( .A(n105), .B(b[22]), .Z(n151) );
  INV_X1 U85 ( .A(a[21]), .ZN(n102) );
  INV_X1 U86 ( .A(b[21]), .ZN(n101) );
  XOR2_X1 U87 ( .A(n102), .B(b[21]), .Z(n149) );
  INV_X1 U88 ( .A(a[20]), .ZN(n100) );
  INV_X1 U89 ( .A(a[19]), .ZN(n98) );
  INV_X1 U90 ( .A(b[19]), .ZN(n97) );
  XOR2_X1 U91 ( .A(n98), .B(b[19]), .Z(n146) );
  INV_X1 U92 ( .A(a[18]), .ZN(n96) );
  INV_X1 U93 ( .A(b[18]), .ZN(n95) );
  INV_X1 U94 ( .A(a[17]), .ZN(n94) );
  INV_X1 U95 ( .A(b[17]), .ZN(n93) );
  XOR2_X1 U96 ( .A(n94), .B(b[17]), .Z(n142) );
  INV_X1 U97 ( .A(a[16]), .ZN(n91) );
  INV_X1 U98 ( .A(b[16]), .ZN(n90) );
  XOR2_X1 U99 ( .A(n91), .B(b[16]), .Z(n141) );
  INV_X1 U100 ( .A(a[15]), .ZN(n89) );
  INV_X1 U101 ( .A(b[15]), .ZN(n88) );
  INV_X1 U102 ( .A(a[14]), .ZN(n87) );
  INV_X1 U103 ( .A(b[14]), .ZN(n86) );
  XOR2_X1 U104 ( .A(n87), .B(b[14]), .Z(n138) );
  INV_X1 U105 ( .A(a[13]), .ZN(n85) );
  INV_X1 U106 ( .A(b[13]), .ZN(n84) );
  INV_X1 U107 ( .A(a[12]), .ZN(n83) );
  INV_X1 U108 ( .A(b[12]), .ZN(n82) );
  XOR2_X1 U109 ( .A(n83), .B(b[12]), .Z(n135) );
  INV_X1 U110 ( .A(a[11]), .ZN(n81) );
  INV_X1 U111 ( .A(b[11]), .ZN(n80) );
  XOR2_X1 U112 ( .A(n81), .B(b[11]), .Z(n133) );
  INV_X1 U113 ( .A(a[10]), .ZN(n78) );
  INV_X1 U114 ( .A(b[10]), .ZN(n77) );
  XOR2_X1 U115 ( .A(n78), .B(b[10]), .Z(n132) );
  INV_X1 U116 ( .A(a[9]), .ZN(n76) );
  INV_X1 U117 ( .A(b[9]), .ZN(n75) );
  INV_X1 U118 ( .A(a[8]), .ZN(n74) );
  INV_X1 U119 ( .A(b[8]), .ZN(n73) );
  XOR2_X1 U120 ( .A(n74), .B(b[8]), .Z(n128) );
  INV_X1 U121 ( .A(a[7]), .ZN(n71) );
  INV_X1 U122 ( .A(b[7]), .ZN(n70) );
  XOR2_X1 U123 ( .A(n71), .B(b[7]), .Z(n126) );
  INV_X1 U124 ( .A(a[6]), .ZN(n68) );
  INV_X1 U125 ( .A(b[6]), .ZN(n67) );
  XOR2_X1 U126 ( .A(n68), .B(b[6]), .Z(n124) );
  INV_X1 U127 ( .A(a[5]), .ZN(n65) );
  INV_X1 U128 ( .A(b[5]), .ZN(n64) );
  XOR2_X1 U129 ( .A(n65), .B(b[5]), .Z(n122) );
  INV_X1 U130 ( .A(a[4]), .ZN(n62) );
  INV_X1 U131 ( .A(b[4]), .ZN(n61) );
  XOR2_X1 U132 ( .A(n62), .B(b[4]), .Z(n119) );
  INV_X1 U133 ( .A(a[3]), .ZN(n59) );
  INV_X1 U134 ( .A(b[3]), .ZN(n58) );
  XOR2_X1 U135 ( .A(n59), .B(b[3]), .Z(n116) );
  INV_X1 U136 ( .A(a[2]), .ZN(n56) );
  INV_X1 U137 ( .A(b[2]), .ZN(n55) );
  INV_X1 U138 ( .A(a[1]), .ZN(n54) );
  INV_X1 U139 ( .A(b[1]), .ZN(n53) );
  INV_X1 U140 ( .A(a[0]), .ZN(n51) );
  INV_X1 U141 ( .A(b[0]), .ZN(n50) );
  XOR2_X1 U142 ( .A(b[0]), .B(n51), .Z(n109) );
  INV_X1 U143 ( .A(cin), .ZN(n49) );
  OAI22_X1 U144 ( .A1(n51), .A2(n50), .B1(n109), .B2(n49), .ZN(n112) );
  INV_X1 U145 ( .A(n112), .ZN(n52) );
  OAI22_X1 U146 ( .A1(n53), .A2(n54), .B1(n110), .B2(n52), .ZN(n115) );
  OAI22_X1 U147 ( .A1(n56), .A2(n55), .B1(n18), .B2(n113), .ZN(n118) );
  INV_X1 U148 ( .A(n118), .ZN(n57) );
  OAI22_X1 U149 ( .A1(n59), .A2(n58), .B1(n57), .B2(n116), .ZN(n121) );
  INV_X1 U150 ( .A(n121), .ZN(n60) );
  OAI22_X1 U151 ( .A1(n62), .A2(n61), .B1(n60), .B2(n119), .ZN(n123) );
  INV_X1 U152 ( .A(n123), .ZN(n63) );
  OAI22_X1 U153 ( .A1(n65), .A2(n64), .B1(n63), .B2(n122), .ZN(n125) );
  INV_X1 U154 ( .A(n125), .ZN(n66) );
  OAI22_X1 U155 ( .A1(n68), .A2(n67), .B1(n66), .B2(n124), .ZN(n127) );
  INV_X1 U156 ( .A(n127), .ZN(n69) );
  OAI22_X1 U157 ( .A1(n71), .A2(n70), .B1(n69), .B2(n126), .ZN(n129) );
  INV_X1 U158 ( .A(n129), .ZN(n72) );
  OAI22_X1 U159 ( .A1(n74), .A2(n73), .B1(n72), .B2(n128), .ZN(n131) );
  OAI22_X1 U160 ( .A1(n78), .A2(n77), .B1(n8), .B2(n132), .ZN(n134) );
  INV_X1 U161 ( .A(n134), .ZN(n79) );
  OAI22_X1 U162 ( .A1(n91), .A2(n90), .B1(n14), .B2(n141), .ZN(n143) );
  INV_X1 U163 ( .A(n143), .ZN(n92) );
  OAI22_X1 U164 ( .A1(n94), .A2(n93), .B1(n92), .B2(n142), .ZN(n145) );
  OAI22_X1 U165 ( .A1(n98), .A2(n97), .B1(n15), .B2(n146), .ZN(n148) );
  INV_X1 U166 ( .A(n148), .ZN(n99) );
  OAI22_X1 U167 ( .A1(n105), .A2(n104), .B1(n103), .B2(n151), .ZN(n153) );
  INV_X1 U168 ( .A(n40), .ZN(n108) );
  INV_X1 U169 ( .A(b[23]), .ZN(n106) );
  OAI22_X1 U170 ( .A1(n108), .A2(n152), .B1(n107), .B2(n106), .ZN(cout) );
  INV_X1 U171 ( .A(n110), .ZN(n111) );
  XOR2_X1 U172 ( .A(n112), .B(n111), .Z(result[1]) );
  INV_X1 U173 ( .A(n113), .ZN(n114) );
  XOR2_X1 U174 ( .A(n31), .B(n114), .Z(result[2]) );
  INV_X1 U175 ( .A(n116), .ZN(n117) );
  XOR2_X1 U176 ( .A(n32), .B(n117), .Z(result[3]) );
  INV_X1 U177 ( .A(n119), .ZN(n120) );
  XOR2_X1 U178 ( .A(n26), .B(n120), .Z(result[4]) );
endmodule


module comparator24bit_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n2, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17, n18, n19,
         n20, n21, n23, n24, n25, n26, n27, n28, n30, n31, n32, n33, n35, n37,
         n38, n39, n40, n41, n44, n45, n46, n47, n48, n49, n50, n52, n54, n55,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n160, n161, n162, n163, n164;

  NAND2_X1 U97 ( .A1(n63), .A2(n149), .ZN(n150) );
  NAND2_X1 U98 ( .A1(n148), .A2(n156), .ZN(n151) );
  NAND2_X1 U99 ( .A1(n150), .A2(n151), .ZN(DIFF[5]) );
  INV_X1 U100 ( .A(n63), .ZN(n148) );
  INV_X1 U101 ( .A(n156), .ZN(n149) );
  AND4_X1 U102 ( .A1(n54), .A2(n46), .A3(n38), .A4(n30), .ZN(n28) );
  CLKBUF_X1 U103 ( .A(B[5]), .Z(n156) );
  OR2_X2 U104 ( .A1(n66), .A2(n58), .ZN(n157) );
  NAND2_X1 U105 ( .A1(n28), .A2(n57), .ZN(n152) );
  NAND2_X1 U106 ( .A1(n28), .A2(n57), .ZN(n27) );
  BUF_X1 U107 ( .A(B[8]), .Z(n153) );
  OR2_X1 U108 ( .A1(B[6]), .A2(n154), .ZN(n155) );
  INV_X1 U109 ( .A(n62), .ZN(n154) );
  OR2_X1 U110 ( .A1(n158), .A2(n154), .ZN(n61) );
  BUF_X1 U111 ( .A(n66), .Z(n158) );
  CLKBUF_X1 U112 ( .A(B[0]), .Z(DIFF[0]) );
  NOR2_X1 U113 ( .A1(n66), .A2(n58), .ZN(n57) );
  XNOR2_X1 U114 ( .A(n160), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U115 ( .A1(n157), .A2(n35), .ZN(n160) );
  OR2_X1 U116 ( .A1(B[8]), .A2(B[9]), .ZN(n161) );
  CLKBUF_X1 U117 ( .A(B[4]), .Z(n162) );
  OR2_X1 U118 ( .A1(n16), .A2(n5), .ZN(n163) );
  XOR2_X1 U119 ( .A(n164), .B(n41), .Z(DIFF[12]) );
  NOR2_X1 U120 ( .A1(n157), .A2(n45), .ZN(n164) );
  INV_X1 U121 ( .A(n38), .ZN(n37) );
  INV_X1 U122 ( .A(n45), .ZN(n44) );
  INV_X1 U123 ( .A(n16), .ZN(n15) );
  INV_X1 U124 ( .A(n24), .ZN(n23) );
  INV_X1 U125 ( .A(n25), .ZN(n24) );
  NAND2_X1 U126 ( .A1(n9), .A2(n6), .ZN(n5) );
  INV_X1 U127 ( .A(B[22]), .ZN(n6) );
  INV_X1 U128 ( .A(n161), .ZN(n52) );
  NAND2_X1 U129 ( .A1(n65), .A2(n64), .ZN(n63) );
  INV_X1 U130 ( .A(n162), .ZN(n64) );
  NOR2_X1 U131 ( .A1(B[8]), .A2(B[9]), .ZN(n54) );
  NAND2_X1 U132 ( .A1(n23), .A2(n20), .ZN(n19) );
  INV_X1 U133 ( .A(B[18]), .ZN(n20) );
  NAND2_X1 U134 ( .A1(n15), .A2(n12), .ZN(n11) );
  INV_X1 U135 ( .A(B[20]), .ZN(n12) );
  INV_X1 U136 ( .A(B[10]), .ZN(n49) );
  XOR2_X1 U137 ( .A(n152), .B(B[16]), .Z(DIFF[16]) );
  NOR2_X1 U138 ( .A1(B[16]), .A2(B[17]), .ZN(n25) );
  NOR2_X1 U139 ( .A1(n37), .A2(B[14]), .ZN(n33) );
  NOR2_X1 U140 ( .A1(B[20]), .A2(B[21]), .ZN(n9) );
  INV_X1 U141 ( .A(n158), .ZN(n65) );
  NAND2_X1 U142 ( .A1(n54), .A2(n46), .ZN(n45) );
  NAND2_X1 U143 ( .A1(n25), .A2(n17), .ZN(n16) );
  NOR2_X1 U144 ( .A1(B[18]), .A2(B[19]), .ZN(n17) );
  NOR2_X1 U145 ( .A1(B[14]), .A2(B[15]), .ZN(n30) );
  XNOR2_X1 U146 ( .A(n68), .B(B[3]), .ZN(DIFF[3]) );
  NAND2_X1 U147 ( .A1(n15), .A2(n9), .ZN(n8) );
  INV_X1 U148 ( .A(B[12]), .ZN(n41) );
  NAND2_X1 U149 ( .A1(n44), .A2(n41), .ZN(n40) );
  NAND2_X1 U150 ( .A1(n44), .A2(n38), .ZN(n35) );
  NOR2_X1 U151 ( .A1(n27), .A2(n163), .ZN(n2) );
  XNOR2_X1 U152 ( .A(n2), .B(B[23]), .ZN(DIFF[23]) );
  NAND2_X1 U153 ( .A1(n52), .A2(n49), .ZN(n48) );
  XNOR2_X1 U154 ( .A(n39), .B(B[13]), .ZN(DIFF[13]) );
  NOR2_X1 U155 ( .A1(n157), .A2(n40), .ZN(n39) );
  NOR2_X1 U156 ( .A1(n157), .A2(n32), .ZN(n31) );
  NAND2_X1 U157 ( .A1(n33), .A2(n44), .ZN(n32) );
  INV_X1 U158 ( .A(n70), .ZN(n69) );
  XNOR2_X1 U159 ( .A(n31), .B(B[15]), .ZN(DIFF[15]) );
  NOR2_X1 U160 ( .A1(B[1]), .A2(B[0]), .ZN(n70) );
  NOR2_X1 U161 ( .A1(n152), .A2(n8), .ZN(n7) );
  NOR2_X1 U162 ( .A1(n157), .A2(n161), .ZN(n50) );
  XNOR2_X1 U163 ( .A(n60), .B(B[7]), .ZN(DIFF[7]) );
  XNOR2_X1 U164 ( .A(n21), .B(B[18]), .ZN(DIFF[18]) );
  XNOR2_X1 U165 ( .A(n13), .B(B[20]), .ZN(DIFF[20]) );
  XNOR2_X1 U166 ( .A(n26), .B(B[17]), .ZN(DIFF[17]) );
  XOR2_X1 U167 ( .A(n61), .B(B[6]), .Z(DIFF[6]) );
  NOR2_X1 U168 ( .A1(n155), .A2(n158), .ZN(n60) );
  NOR2_X1 U169 ( .A1(B[6]), .A2(B[7]), .ZN(n59) );
  XNOR2_X1 U170 ( .A(n55), .B(B[9]), .ZN(DIFF[9]) );
  XNOR2_X1 U171 ( .A(n50), .B(B[10]), .ZN(DIFF[10]) );
  XNOR2_X1 U172 ( .A(n18), .B(B[19]), .ZN(DIFF[19]) );
  NOR2_X1 U173 ( .A1(B[10]), .A2(B[11]), .ZN(n46) );
  XNOR2_X1 U174 ( .A(n10), .B(B[21]), .ZN(DIFF[21]) );
  NOR2_X1 U175 ( .A1(B[12]), .A2(B[13]), .ZN(n38) );
  XNOR2_X1 U176 ( .A(n47), .B(B[11]), .ZN(DIFF[11]) );
  NOR2_X1 U177 ( .A1(n157), .A2(n48), .ZN(n47) );
  NOR2_X1 U178 ( .A1(n27), .A2(n11), .ZN(n10) );
  NOR2_X1 U179 ( .A1(n27), .A2(n19), .ZN(n18) );
  NOR2_X1 U180 ( .A1(n152), .A2(B[16]), .ZN(n26) );
  NOR2_X1 U181 ( .A1(n152), .A2(n16), .ZN(n13) );
  NOR2_X1 U182 ( .A1(n152), .A2(n24), .ZN(n21) );
  XNOR2_X1 U183 ( .A(n7), .B(B[22]), .ZN(DIFF[22]) );
  XOR2_X1 U184 ( .A(n157), .B(n153), .Z(DIFF[8]) );
  NOR2_X1 U185 ( .A1(n157), .A2(n153), .ZN(n55) );
  XNOR2_X1 U186 ( .A(n65), .B(n162), .ZN(DIFF[4]) );
  NAND2_X1 U187 ( .A1(n62), .A2(n59), .ZN(n58) );
  NOR2_X1 U188 ( .A1(B[4]), .A2(B[5]), .ZN(n62) );
  NOR2_X1 U189 ( .A1(B[2]), .A2(B[3]), .ZN(n67) );
  XOR2_X1 U190 ( .A(n69), .B(B[2]), .Z(DIFF[2]) );
  NOR2_X1 U191 ( .A1(n69), .A2(B[2]), .ZN(n68) );
  NAND2_X1 U192 ( .A1(n67), .A2(n70), .ZN(n66) );
  XOR2_X1 U193 ( .A(B[1]), .B(DIFF[0]), .Z(DIFF[1]) );
endmodule


module comparator24bit_DW01_add_1 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;
  wire   n1, n4, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n24, n25, n26, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n148,
         n149, n150, n151;

  OAI22_X1 U95 ( .A1(A[18]), .A2(B[18]), .B1(A[19]), .B2(B[19]), .ZN(n148) );
  INV_X1 U96 ( .A(n148), .ZN(n150) );
  OAI22_X1 U97 ( .A1(A[22]), .A2(B[22]), .B1(A[23]), .B2(B[23]), .ZN(n149) );
  INV_X1 U98 ( .A(n149), .ZN(n9) );
  AOI21_X1 U99 ( .B1(n81), .B2(n87), .A(n82), .ZN(n80) );
  NOR2_X1 U100 ( .A1(A[5]), .A2(B[5]), .ZN(n76) );
  NOR2_X1 U101 ( .A1(A[3]), .A2(B[3]), .ZN(n83) );
  NAND2_X1 U102 ( .A1(A[4]), .A2(B[4]), .ZN(n79) );
  NAND2_X1 U103 ( .A1(A[5]), .A2(B[5]), .ZN(n77) );
  NAND2_X1 U104 ( .A1(A[8]), .A2(B[8]), .ZN(n64) );
  NAND2_X1 U105 ( .A1(A[6]), .A2(B[6]), .ZN(n73) );
  NAND2_X1 U106 ( .A1(B[7]), .A2(A[7]), .ZN(n71) );
  OAI21_X1 U107 ( .B1(n88), .B2(n90), .A(n89), .ZN(n87) );
  NAND2_X1 U108 ( .A1(A[1]), .A2(B[1]), .ZN(n89) );
  NOR2_X1 U109 ( .A1(A[1]), .A2(B[1]), .ZN(n88) );
  OAI21_X1 U110 ( .B1(n83), .B2(n86), .A(n84), .ZN(n82) );
  NAND2_X1 U111 ( .A1(A[2]), .A2(B[2]), .ZN(n86) );
  NAND2_X1 U112 ( .A1(A[3]), .A2(B[3]), .ZN(n84) );
  NOR2_X1 U113 ( .A1(n70), .A2(n72), .ZN(n68) );
  NOR2_X1 U114 ( .A1(A[6]), .A2(B[6]), .ZN(n72) );
  NOR2_X1 U115 ( .A1(A[8]), .A2(B[8]), .ZN(n63) );
  NOR2_X1 U116 ( .A1(n85), .A2(n83), .ZN(n81) );
  NOR2_X1 U117 ( .A1(A[2]), .A2(B[2]), .ZN(n85) );
  NOR2_X1 U118 ( .A1(n78), .A2(n76), .ZN(n74) );
  NOR2_X1 U119 ( .A1(A[4]), .A2(B[4]), .ZN(n78) );
  OR2_X1 U120 ( .A1(n7), .A2(n21), .ZN(n151) );
  NAND2_X1 U121 ( .A1(A[16]), .A2(B[16]), .ZN(n34) );
  NOR2_X1 U122 ( .A1(A[16]), .A2(B[16]), .ZN(n33) );
  OAI21_X1 U123 ( .B1(n31), .B2(n34), .A(n32), .ZN(n30) );
  OAI21_X1 U124 ( .B1(n17), .B2(n20), .A(n18), .ZN(n16) );
  NOR2_X1 U125 ( .A1(A[21]), .A2(B[21]), .ZN(n17) );
  NAND2_X1 U126 ( .A1(n59), .A2(n53), .ZN(n51) );
  NOR2_X1 U127 ( .A1(n57), .A2(n55), .ZN(n53) );
  NAND2_X1 U128 ( .A1(A[10]), .A2(B[10]), .ZN(n58) );
  AOI21_X1 U129 ( .B1(n150), .B2(n30), .A(n24), .ZN(n22) );
  NAND2_X1 U130 ( .A1(A[13]), .A2(B[13]), .ZN(n48) );
  NAND2_X1 U131 ( .A1(A[20]), .A2(B[20]), .ZN(n20) );
  NAND2_X1 U132 ( .A1(A[14]), .A2(B[14]), .ZN(n44) );
  NAND2_X1 U133 ( .A1(A[11]), .A2(B[11]), .ZN(n56) );
  NAND2_X1 U134 ( .A1(A[12]), .A2(B[12]), .ZN(n50) );
  OAI21_X1 U135 ( .B1(n11), .B2(n14), .A(n12), .ZN(n10) );
  OAI21_X1 U136 ( .B1(n80), .B2(n66), .A(n67), .ZN(n65) );
  NAND2_X1 U137 ( .A1(n68), .A2(n74), .ZN(n66) );
  AOI21_X1 U138 ( .B1(n68), .B2(n75), .A(n69), .ZN(n67) );
  OAI21_X1 U139 ( .B1(n76), .B2(n79), .A(n77), .ZN(n75) );
  OAI21_X1 U140 ( .B1(n70), .B2(n73), .A(n71), .ZN(n69) );
  NOR2_X1 U141 ( .A1(A[13]), .A2(B[13]), .ZN(n47) );
  NOR2_X1 U142 ( .A1(A[12]), .A2(B[12]), .ZN(n49) );
  OAI21_X1 U143 ( .B1(n41), .B2(n44), .A(n42), .ZN(n40) );
  OAI21_X1 U144 ( .B1(n55), .B2(n58), .A(n56), .ZN(n54) );
  NOR2_X1 U145 ( .A1(B[7]), .A2(A[7]), .ZN(n70) );
  OAI21_X1 U146 ( .B1(n61), .B2(n64), .A(n62), .ZN(n60) );
  NOR2_X1 U147 ( .A1(n63), .A2(n61), .ZN(n59) );
  NAND2_X1 U148 ( .A1(A[9]), .A2(B[9]), .ZN(n62) );
  NOR2_X1 U149 ( .A1(A[9]), .A2(B[9]), .ZN(n61) );
  OAI21_X1 U150 ( .B1(n22), .B2(n7), .A(n8), .ZN(n6) );
  NAND2_X1 U151 ( .A1(n9), .A2(n15), .ZN(n7) );
  OAI21_X1 U152 ( .B1(n25), .B2(n28), .A(n26), .ZN(n24) );
  NAND2_X1 U153 ( .A1(A[18]), .A2(B[18]), .ZN(n28) );
  NOR2_X1 U154 ( .A1(A[20]), .A2(B[20]), .ZN(n19) );
  NOR2_X1 U155 ( .A1(n19), .A2(n17), .ZN(n15) );
  NOR2_X1 U156 ( .A1(n33), .A2(n31), .ZN(n29) );
  NAND2_X1 U157 ( .A1(A[17]), .A2(B[17]), .ZN(n32) );
  NOR2_X1 U158 ( .A1(A[17]), .A2(B[17]), .ZN(n31) );
  NOR2_X1 U159 ( .A1(n51), .A2(n37), .ZN(n35) );
  OAI21_X1 U160 ( .B1(n52), .B2(n37), .A(n38), .ZN(n36) );
  AOI21_X1 U161 ( .B1(n9), .B2(n16), .A(n10), .ZN(n8) );
  NAND2_X1 U162 ( .A1(A[23]), .A2(B[23]), .ZN(n12) );
  NOR2_X1 U163 ( .A1(A[23]), .A2(B[23]), .ZN(n11) );
  NOR2_X1 U164 ( .A1(A[10]), .A2(B[10]), .ZN(n57) );
  AOI21_X1 U165 ( .B1(n65), .B2(n35), .A(n36), .ZN(n1) );
  INV_X1 U166 ( .A(n6), .ZN(n4) );
  NAND2_X1 U167 ( .A1(A[19]), .A2(B[19]), .ZN(n26) );
  NOR2_X1 U168 ( .A1(A[19]), .A2(B[19]), .ZN(n25) );
  OAI21_X1 U169 ( .B1(n1), .B2(n151), .A(n4), .ZN(SUM[24]) );
  AOI21_X1 U170 ( .B1(n39), .B2(n46), .A(n40), .ZN(n38) );
  NAND2_X1 U171 ( .A1(n45), .A2(n39), .ZN(n37) );
  NAND2_X1 U172 ( .A1(A[21]), .A2(B[21]), .ZN(n18) );
  AOI21_X1 U173 ( .B1(n53), .B2(n60), .A(n54), .ZN(n52) );
  NOR2_X1 U174 ( .A1(A[11]), .A2(B[11]), .ZN(n55) );
  OAI21_X1 U175 ( .B1(n47), .B2(n50), .A(n48), .ZN(n46) );
  NOR2_X1 U176 ( .A1(n49), .A2(n47), .ZN(n45) );
  NOR2_X1 U177 ( .A1(n41), .A2(n43), .ZN(n39) );
  NOR2_X1 U178 ( .A1(A[14]), .A2(B[14]), .ZN(n43) );
  NAND2_X1 U179 ( .A1(A[15]), .A2(B[15]), .ZN(n42) );
  NOR2_X1 U180 ( .A1(B[15]), .A2(A[15]), .ZN(n41) );
  NAND2_X1 U181 ( .A1(A[22]), .A2(B[22]), .ZN(n14) );
  NAND2_X1 U182 ( .A1(n29), .A2(n150), .ZN(n21) );
  NAND2_X1 U183 ( .A1(A[0]), .A2(B[0]), .ZN(n90) );
endmodule


module comparator24bit ( a, b, f_bigger );
  input [23:0] a;
  input [23:0] b;
  output f_bigger;
  wire   complement_b_9_, complement_b_8_, complement_b_7_, complement_b_6_,
         complement_b_5_, complement_b_4_, complement_b_3_, complement_b_2_,
         complement_b_23_, complement_b_22_, complement_b_21_,
         complement_b_20_, complement_b_1_, complement_b_19_, complement_b_18_,
         complement_b_17_, complement_b_16_, complement_b_15_,
         complement_b_14_, complement_b_13_, complement_b_12_,
         complement_b_11_, complement_b_10_, complement_b_0_,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24;

  comparator24bit_DW01_sub_1 sub_add_11_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(b), .CI(1'b0), .DIFF({
        complement_b_23_, complement_b_22_, complement_b_21_, complement_b_20_, 
        complement_b_19_, complement_b_18_, complement_b_17_, complement_b_16_, 
        complement_b_15_, complement_b_14_, complement_b_13_, complement_b_12_, 
        complement_b_11_, complement_b_10_, complement_b_9_, complement_b_8_, 
        complement_b_7_, complement_b_6_, complement_b_5_, complement_b_4_, 
        complement_b_3_, complement_b_2_, complement_b_1_, complement_b_0_})
         );
  comparator24bit_DW01_add_1 add_13 ( .A({1'b0, a}), .B({1'b0, 
        complement_b_23_, complement_b_22_, complement_b_21_, complement_b_20_, 
        complement_b_19_, complement_b_18_, complement_b_17_, complement_b_16_, 
        complement_b_15_, complement_b_14_, complement_b_13_, complement_b_12_, 
        complement_b_11_, complement_b_10_, complement_b_9_, complement_b_8_, 
        complement_b_7_, complement_b_6_, complement_b_5_, complement_b_4_, 
        complement_b_3_, complement_b_2_, complement_b_1_, complement_b_0_}), 
        .CI(1'b0), .SUM({f_bigger, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24}) );
endmodule


module Adder24Bit_DW01_add_5 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n25, n106, n107, n108, n110, n111;

  HA_X1 U2 ( .A(n3), .B(A[22]), .CO(n2), .S(SUM[22]) );
  HA_X1 U3 ( .A(n4), .B(A[21]), .CO(n3), .S(SUM[21]) );
  HA_X1 U4 ( .A(n5), .B(A[20]), .CO(n4), .S(SUM[20]) );
  HA_X1 U5 ( .A(n6), .B(A[19]), .CO(n5), .S(SUM[19]) );
  HA_X1 U7 ( .A(n8), .B(A[17]), .CO(n7), .S(SUM[17]) );
  HA_X1 U8 ( .A(n9), .B(A[16]), .CO(n8), .S(SUM[16]) );
  HA_X1 U9 ( .A(n10), .B(A[15]), .CO(n9), .S(SUM[15]) );
  HA_X1 U12 ( .A(n13), .B(A[12]), .CO(n12), .S(SUM[12]) );
  HA_X1 U13 ( .A(n14), .B(A[11]), .CO(n13), .S(SUM[11]) );
  HA_X1 U14 ( .A(n15), .B(A[10]), .CO(n14), .S(SUM[10]) );
  HA_X1 U15 ( .A(n16), .B(A[9]), .CO(n15), .S(SUM[9]) );
  HA_X1 U16 ( .A(n17), .B(A[8]), .CO(n16), .S(SUM[8]) );
  HA_X1 U17 ( .A(n18), .B(A[7]), .CO(n17), .S(SUM[7]) );
  HA_X1 U18 ( .A(n19), .B(A[6]), .CO(n18), .S(SUM[6]) );
  HA_X1 U19 ( .A(n20), .B(A[5]), .CO(n19), .S(SUM[5]) );
  HA_X1 U20 ( .A(n21), .B(A[4]), .CO(n20), .S(SUM[4]) );
  HA_X1 U21 ( .A(n22), .B(A[3]), .CO(n21), .S(SUM[3]) );
  HA_X1 U22 ( .A(n108), .B(A[2]), .CO(n22), .S(SUM[2]) );
  XOR2_X1 U33 ( .A(n12), .B(A[13]), .Z(SUM[13]) );
  INV_X1 U34 ( .A(n106), .ZN(n11) );
  NAND2_X1 U35 ( .A1(n12), .A2(A[13]), .ZN(n106) );
  XOR2_X1 U36 ( .A(n11), .B(A[14]), .Z(SUM[14]) );
  XOR2_X1 U37 ( .A(n7), .B(A[18]), .Z(SUM[18]) );
  INV_X1 U38 ( .A(n107), .ZN(n6) );
  NAND2_X1 U39 ( .A1(n7), .A2(A[18]), .ZN(n107) );
  AND2_X1 U40 ( .A1(n110), .A2(A[1]), .ZN(n108) );
  AND2_X1 U41 ( .A1(n11), .A2(A[14]), .ZN(n10) );
  XOR2_X1 U42 ( .A(n110), .B(A[1]), .Z(SUM[1]) );
  AND2_X1 U43 ( .A1(n25), .A2(n111), .ZN(SUM[0]) );
  AND2_X1 U44 ( .A1(A[0]), .A2(B[0]), .ZN(n110) );
  XOR2_X1 U45 ( .A(n2), .B(A[23]), .Z(SUM[23]) );
  OR2_X1 U46 ( .A1(A[0]), .A2(B[0]), .ZN(n111) );
  NAND2_X1 U47 ( .A1(A[0]), .A2(B[0]), .ZN(n25) );
endmodule


module Adder24Bit_DW01_add_4 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;
  wire   n3, n5, n6, n7, n8, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n116, n117,
         n118, n119, n120, n121, n123;

  HA_X1 U15 ( .A(n13), .B(A[19]), .CO(n12), .S(SUM[19]) );
  HA_X1 U16 ( .A(n14), .B(A[18]), .S(SUM[18]) );
  HA_X1 U17 ( .A(n15), .B(A[17]), .CO(n14), .S(SUM[17]) );
  HA_X1 U18 ( .A(n16), .B(A[16]), .CO(n15), .S(SUM[16]) );
  HA_X1 U19 ( .A(n17), .B(A[15]), .S(SUM[15]) );
  HA_X1 U20 ( .A(n18), .B(A[14]), .CO(n17), .S(SUM[14]) );
  HA_X1 U21 ( .A(n19), .B(A[13]), .CO(n18), .S(SUM[13]) );
  HA_X1 U22 ( .A(A[12]), .B(n20), .CO(n19), .S(SUM[12]) );
  HA_X1 U23 ( .A(A[11]), .B(n21), .CO(n20), .S(SUM[11]) );
  HA_X1 U24 ( .A(n22), .B(A[10]), .CO(n21), .S(SUM[10]) );
  HA_X1 U25 ( .A(n23), .B(A[9]), .CO(n22), .S(SUM[9]) );
  HA_X1 U26 ( .A(n24), .B(A[8]), .CO(n23), .S(SUM[8]) );
  HA_X1 U27 ( .A(n25), .B(A[7]), .CO(n24), .S(SUM[7]) );
  HA_X1 U28 ( .A(n26), .B(A[6]), .CO(n25), .S(SUM[6]) );
  HA_X1 U29 ( .A(n27), .B(A[5]), .CO(n26), .S(SUM[5]) );
  HA_X1 U30 ( .A(n28), .B(A[4]), .CO(n27), .S(SUM[4]) );
  HA_X1 U31 ( .A(n29), .B(A[3]), .CO(n28), .S(SUM[3]) );
  HA_X1 U32 ( .A(n30), .B(A[2]), .CO(n29), .S(SUM[2]) );
  HA_X1 U33 ( .A(n31), .B(A[1]), .CO(n30), .S(SUM[1]) );
  AND3_X1 U43 ( .A1(A[18]), .A2(A[17]), .A3(A[16]), .ZN(n116) );
  AND2_X2 U44 ( .A1(n16), .A2(n116), .ZN(n13) );
  AND3_X2 U45 ( .A1(n18), .A2(A[14]), .A3(A[15]), .ZN(n16) );
  AND3_X1 U46 ( .A1(A[22]), .A2(n120), .A3(n12), .ZN(n6) );
  CLKBUF_X1 U47 ( .A(n6), .Z(n117) );
  AND2_X1 U48 ( .A1(n13), .A2(A[19]), .ZN(n118) );
  AND2_X1 U49 ( .A1(n13), .A2(A[19]), .ZN(n119) );
  AND2_X1 U50 ( .A1(A[20]), .A2(A[21]), .ZN(n120) );
  XOR2_X1 U51 ( .A(A[20]), .B(n119), .Z(SUM[20]) );
  AND2_X1 U52 ( .A1(A[20]), .A2(n118), .ZN(n121) );
  INV_X1 U53 ( .A(A[22]), .ZN(n7) );
  XNOR2_X1 U54 ( .A(n3), .B(A[24]), .ZN(SUM[24]) );
  AND2_X1 U55 ( .A1(n123), .A2(n33), .ZN(SUM[0]) );
  XOR2_X1 U56 ( .A(A[21]), .B(n121), .Z(SUM[21]) );
  OR2_X1 U57 ( .A1(A[0]), .A2(B[0]), .ZN(n123) );
  XNOR2_X1 U58 ( .A(n5), .B(n117), .ZN(SUM[23]) );
  INV_X1 U59 ( .A(A[23]), .ZN(n5) );
  NAND2_X1 U60 ( .A1(A[23]), .A2(n6), .ZN(n3) );
  XOR2_X1 U61 ( .A(n7), .B(n8), .Z(SUM[22]) );
  INV_X1 U62 ( .A(n33), .ZN(n31) );
  NAND2_X1 U63 ( .A1(A[0]), .A2(B[0]), .ZN(n33) );
  NAND2_X1 U64 ( .A1(n120), .A2(n12), .ZN(n8) );
endmodule


module Adder24Bit_DW01_add_6 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n25, n26, n106;

  HA_X1 U2 ( .A(n3), .B(A[22]), .CO(n2), .S(SUM[22]) );
  HA_X1 U3 ( .A(n4), .B(A[21]), .CO(n3), .S(SUM[21]) );
  HA_X1 U4 ( .A(n5), .B(A[20]), .CO(n4), .S(SUM[20]) );
  HA_X1 U5 ( .A(n6), .B(A[19]), .CO(n5), .S(SUM[19]) );
  HA_X1 U6 ( .A(n7), .B(A[18]), .CO(n6), .S(SUM[18]) );
  HA_X1 U7 ( .A(n8), .B(A[17]), .CO(n7), .S(SUM[17]) );
  HA_X1 U8 ( .A(n9), .B(A[16]), .CO(n8), .S(SUM[16]) );
  HA_X1 U9 ( .A(n10), .B(A[15]), .CO(n9), .S(SUM[15]) );
  HA_X1 U10 ( .A(n11), .B(A[14]), .CO(n10), .S(SUM[14]) );
  HA_X1 U11 ( .A(n12), .B(A[13]), .CO(n11), .S(SUM[13]) );
  HA_X1 U12 ( .A(n13), .B(A[12]), .CO(n12), .S(SUM[12]) );
  HA_X1 U13 ( .A(n14), .B(A[11]), .CO(n13), .S(SUM[11]) );
  HA_X1 U14 ( .A(n15), .B(A[10]), .CO(n14), .S(SUM[10]) );
  HA_X1 U15 ( .A(n16), .B(A[9]), .CO(n15), .S(SUM[9]) );
  HA_X1 U16 ( .A(n17), .B(A[8]), .CO(n16), .S(SUM[8]) );
  HA_X1 U17 ( .A(n18), .B(A[7]), .CO(n17), .S(SUM[7]) );
  HA_X1 U18 ( .A(n19), .B(A[6]), .CO(n18), .S(SUM[6]) );
  HA_X1 U19 ( .A(n20), .B(A[5]), .CO(n19), .S(SUM[5]) );
  HA_X1 U20 ( .A(n21), .B(A[4]), .CO(n20), .S(SUM[4]) );
  HA_X1 U21 ( .A(n22), .B(A[3]), .CO(n21), .S(SUM[3]) );
  HA_X1 U22 ( .A(n23), .B(A[2]), .CO(n22), .S(SUM[2]) );
  HA_X1 U23 ( .A(n26), .B(A[1]), .CO(n23), .S(SUM[1]) );
  OR2_X1 U33 ( .A1(A[0]), .A2(B[0]), .ZN(n106) );
  AND2_X1 U34 ( .A1(n106), .A2(n25), .ZN(SUM[0]) );
  NAND2_X1 U35 ( .A1(A[0]), .A2(B[0]), .ZN(n25) );
  INV_X1 U36 ( .A(n25), .ZN(n26) );
  XOR2_X1 U37 ( .A(n2), .B(A[23]), .Z(SUM[23]) );
endmodule


module Adder24Bit ( a, b, signFO, signSO, result, finalSign, cout );
  input [23:0] a;
  input [23:0] b;
  output [23:0] result;
  input signFO, signSO;
  output finalSign, cout;
  wire   tempCout, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14,
         N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42,
         N43, N44, N45, N46, N47, N48, N49, f_bigger, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N74, N75, tempResult_adjusted_24_,
         tempResult_adjusted_9_, tempResult_adjusted_8_,
         tempResult_adjusted_7_, tempResult_adjusted_6_,
         tempResult_adjusted_5_, tempResult_adjusted_4_,
         tempResult_adjusted_3_, tempResult_adjusted_2_,
         tempResult_adjusted_23_, tempResult_adjusted_22_,
         tempResult_adjusted_21_, tempResult_adjusted_20_,
         tempResult_adjusted_1_, tempResult_adjusted_19_,
         tempResult_adjusted_18_, tempResult_adjusted_17_,
         tempResult_adjusted_16_, tempResult_adjusted_15_,
         tempResult_adjusted_14_, tempResult_adjusted_13_,
         tempResult_adjusted_12_, tempResult_adjusted_11_,
         tempResult_adjusted_10_, tempResult_adjusted_0_, n1, n2, n3, n4, n6,
         n8, n9, n10, n14, n15, n16, n17;
  wire   [23:0] a_op;
  wire   [23:0] b_op;
  wire   [23:0] tempResult;

  carryLookAheadAdder CL ( .a(a_op), .b(b_op), .cin(1'b0), .result(tempResult), 
        .cout(tempCout) );
  comparator24bit Comp ( .a(a), .b(b), .f_bigger(f_bigger) );
  Adder24Bit_DW01_add_5 add_24 ( .A({N26, N27, N28, N29, N30, N31, N32, N33, 
        N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, 
        N48, N49}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, n10}), .CI(1'b0), .SUM(b_op) );
  Adder24Bit_DW01_add_4 add_33 ( .A({N51, N52, N53, N54, N55, N56, N57, N58, 
        N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, 
        N73, N74, N75}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, n9}), .CI(1'b0), .SUM({tempResult_adjusted_24_, 
        tempResult_adjusted_23_, tempResult_adjusted_22_, 
        tempResult_adjusted_21_, tempResult_adjusted_20_, 
        tempResult_adjusted_19_, tempResult_adjusted_18_, 
        tempResult_adjusted_17_, tempResult_adjusted_16_, 
        tempResult_adjusted_15_, tempResult_adjusted_14_, 
        tempResult_adjusted_13_, tempResult_adjusted_12_, 
        tempResult_adjusted_11_, tempResult_adjusted_10_, 
        tempResult_adjusted_9_, tempResult_adjusted_8_, tempResult_adjusted_7_, 
        tempResult_adjusted_6_, tempResult_adjusted_5_, tempResult_adjusted_4_, 
        tempResult_adjusted_3_, tempResult_adjusted_2_, tempResult_adjusted_1_, 
        tempResult_adjusted_0_}) );
  Adder24Bit_DW01_add_6 add_23 ( .A({N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, 
        N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        signFO}), .CI(1'b0), .SUM(a_op) );
  XOR2_X1 U2 ( .A(b[13]), .B(signSO), .Z(N36) );
  XOR2_X1 U3 ( .A(b[18]), .B(signSO), .Z(N31) );
  XOR2_X1 U4 ( .A(tempResult[20]), .B(finalSign), .Z(N55) );
  BUF_X2 U5 ( .A(n3), .Z(n9) );
  AND2_X2 U6 ( .A1(tempResult_adjusted_24_), .A2(n17), .ZN(cout) );
  CLKBUF_X1 U10 ( .A(n9), .Z(n1) );
  INV_X1 U11 ( .A(finalSign), .ZN(n2) );
  XNOR2_X1 U12 ( .A(tempResult[23]), .B(n2), .ZN(N52) );
  XNOR2_X1 U13 ( .A(b[1]), .B(n14), .ZN(N48) );
  XNOR2_X1 U14 ( .A(n4), .B(finalSign), .ZN(N51) );
  MUX2_X1 U15 ( .A(signSO), .B(signFO), .S(f_bigger), .Z(n3) );
  INV_X2 U16 ( .A(n14), .ZN(n10) );
  XNOR2_X1 U17 ( .A(b[0]), .B(n14), .ZN(N49) );
  NAND2_X1 U18 ( .A1(tempCout), .A2(n17), .ZN(n4) );
  XOR2_X1 U19 ( .A(tempResult[4]), .B(finalSign), .Z(N71) );
  XOR2_X1 U20 ( .A(tempResult[3]), .B(n1), .Z(N72) );
  XOR2_X1 U21 ( .A(tempResult[2]), .B(n1), .Z(N73) );
  OR2_X1 U22 ( .A1(tempResult_adjusted_23_), .A2(n6), .ZN(result[23]) );
  INV_X1 U23 ( .A(n16), .ZN(n15) );
  INV_X1 U24 ( .A(signSO), .ZN(n14) );
  CLKBUF_X1 U25 ( .A(cout), .Z(n6) );
  CLKBUF_X1 U26 ( .A(n6), .Z(n8) );
  BUF_X4 U27 ( .A(n9), .Z(finalSign) );
  INV_X1 U28 ( .A(signFO), .ZN(n16) );
  XOR2_X1 U29 ( .A(signSO), .B(b[23]), .Z(N26) );
  XOR2_X1 U30 ( .A(b[22]), .B(signSO), .Z(N27) );
  XOR2_X1 U31 ( .A(b[21]), .B(signSO), .Z(N28) );
  XOR2_X1 U32 ( .A(b[20]), .B(signSO), .Z(N29) );
  XOR2_X1 U33 ( .A(b[19]), .B(signSO), .Z(N30) );
  XOR2_X1 U34 ( .A(b[17]), .B(signSO), .Z(N32) );
  XOR2_X1 U35 ( .A(b[16]), .B(signSO), .Z(N33) );
  XOR2_X1 U36 ( .A(b[15]), .B(signSO), .Z(N34) );
  XOR2_X1 U37 ( .A(b[14]), .B(signSO), .Z(N35) );
  XOR2_X1 U38 ( .A(b[12]), .B(signSO), .Z(N37) );
  XOR2_X1 U39 ( .A(b[11]), .B(n10), .Z(N38) );
  XOR2_X1 U40 ( .A(b[10]), .B(n10), .Z(N39) );
  XOR2_X1 U41 ( .A(b[9]), .B(n10), .Z(N40) );
  XOR2_X1 U42 ( .A(b[8]), .B(n10), .Z(N41) );
  XOR2_X1 U43 ( .A(b[7]), .B(n10), .Z(N42) );
  XOR2_X1 U44 ( .A(b[6]), .B(n10), .Z(N43) );
  XOR2_X1 U45 ( .A(b[5]), .B(n10), .Z(N44) );
  XOR2_X1 U46 ( .A(b[4]), .B(n10), .Z(N45) );
  XOR2_X1 U47 ( .A(b[3]), .B(n10), .Z(N46) );
  XOR2_X1 U48 ( .A(b[2]), .B(n10), .Z(N47) );
  XOR2_X1 U49 ( .A(n15), .B(a[23]), .Z(N2) );
  XOR2_X1 U50 ( .A(a[22]), .B(n15), .Z(N3) );
  XOR2_X1 U51 ( .A(a[21]), .B(n15), .Z(N4) );
  XOR2_X1 U52 ( .A(a[20]), .B(n15), .Z(N5) );
  XOR2_X1 U53 ( .A(a[19]), .B(n15), .Z(N6) );
  XOR2_X1 U54 ( .A(a[18]), .B(n15), .Z(N7) );
  XOR2_X1 U55 ( .A(a[17]), .B(n15), .Z(N8) );
  XOR2_X1 U56 ( .A(a[16]), .B(n15), .Z(N9) );
  XOR2_X1 U57 ( .A(a[15]), .B(n15), .Z(N10) );
  XOR2_X1 U58 ( .A(a[14]), .B(n15), .Z(N11) );
  XOR2_X1 U59 ( .A(a[13]), .B(n15), .Z(N12) );
  XOR2_X1 U60 ( .A(a[12]), .B(n15), .Z(N13) );
  XOR2_X1 U61 ( .A(a[11]), .B(n15), .Z(N14) );
  XOR2_X1 U62 ( .A(a[10]), .B(n15), .Z(N15) );
  XOR2_X1 U63 ( .A(a[9]), .B(signFO), .Z(N16) );
  XOR2_X1 U64 ( .A(a[8]), .B(signFO), .Z(N17) );
  XOR2_X1 U65 ( .A(a[7]), .B(signFO), .Z(N18) );
  XOR2_X1 U66 ( .A(a[6]), .B(n15), .Z(N19) );
  XOR2_X1 U67 ( .A(a[5]), .B(n15), .Z(N20) );
  XOR2_X1 U68 ( .A(a[4]), .B(n15), .Z(N21) );
  XOR2_X1 U69 ( .A(a[3]), .B(n15), .Z(N22) );
  XOR2_X1 U70 ( .A(a[2]), .B(signFO), .Z(N23) );
  XOR2_X1 U71 ( .A(a[1]), .B(signFO), .Z(N24) );
  XOR2_X1 U72 ( .A(a[0]), .B(signFO), .Z(N25) );
  XOR2_X1 U73 ( .A(n14), .B(n15), .Z(n17) );
  XOR2_X1 U74 ( .A(tempResult[22]), .B(finalSign), .Z(N53) );
  XOR2_X1 U75 ( .A(tempResult[21]), .B(finalSign), .Z(N54) );
  XOR2_X1 U76 ( .A(tempResult[19]), .B(finalSign), .Z(N56) );
  XOR2_X1 U77 ( .A(tempResult[18]), .B(finalSign), .Z(N57) );
  XOR2_X1 U78 ( .A(tempResult[17]), .B(finalSign), .Z(N58) );
  XOR2_X1 U79 ( .A(tempResult[16]), .B(finalSign), .Z(N59) );
  XOR2_X1 U80 ( .A(tempResult[15]), .B(finalSign), .Z(N60) );
  XOR2_X1 U81 ( .A(tempResult[14]), .B(finalSign), .Z(N61) );
  XOR2_X1 U82 ( .A(tempResult[13]), .B(finalSign), .Z(N62) );
  XOR2_X1 U83 ( .A(tempResult[12]), .B(finalSign), .Z(N63) );
  XOR2_X1 U84 ( .A(tempResult[11]), .B(finalSign), .Z(N64) );
  XOR2_X1 U85 ( .A(tempResult[10]), .B(finalSign), .Z(N65) );
  XOR2_X1 U86 ( .A(tempResult[9]), .B(finalSign), .Z(N66) );
  XOR2_X1 U87 ( .A(tempResult[8]), .B(finalSign), .Z(N67) );
  XOR2_X1 U88 ( .A(tempResult[7]), .B(finalSign), .Z(N68) );
  XOR2_X1 U89 ( .A(tempResult[6]), .B(finalSign), .Z(N69) );
  XOR2_X1 U90 ( .A(tempResult[5]), .B(finalSign), .Z(N70) );
  XOR2_X1 U91 ( .A(tempResult[1]), .B(n9), .Z(N74) );
  XOR2_X1 U92 ( .A(tempResult[0]), .B(n3), .Z(N75) );
  MUX2_X1 U93 ( .A(tempResult_adjusted_0_), .B(tempResult_adjusted_1_), .S(n8), 
        .Z(result[0]) );
  MUX2_X1 U94 ( .A(tempResult_adjusted_1_), .B(tempResult_adjusted_2_), .S(n8), 
        .Z(result[1]) );
  MUX2_X1 U95 ( .A(tempResult_adjusted_2_), .B(tempResult_adjusted_3_), .S(n8), 
        .Z(result[2]) );
  MUX2_X1 U96 ( .A(tempResult_adjusted_3_), .B(tempResult_adjusted_4_), .S(n8), 
        .Z(result[3]) );
  MUX2_X1 U97 ( .A(tempResult_adjusted_4_), .B(tempResult_adjusted_5_), .S(n8), 
        .Z(result[4]) );
  MUX2_X1 U98 ( .A(tempResult_adjusted_5_), .B(tempResult_adjusted_6_), .S(n8), 
        .Z(result[5]) );
  MUX2_X1 U99 ( .A(tempResult_adjusted_6_), .B(tempResult_adjusted_7_), .S(n8), 
        .Z(result[6]) );
  MUX2_X1 U100 ( .A(tempResult_adjusted_7_), .B(tempResult_adjusted_8_), .S(n8), .Z(result[7]) );
  MUX2_X1 U101 ( .A(tempResult_adjusted_8_), .B(tempResult_adjusted_9_), .S(n8), .Z(result[8]) );
  MUX2_X1 U102 ( .A(tempResult_adjusted_9_), .B(tempResult_adjusted_10_), .S(
        n8), .Z(result[9]) );
  MUX2_X1 U103 ( .A(tempResult_adjusted_10_), .B(tempResult_adjusted_11_), .S(
        n8), .Z(result[10]) );
  MUX2_X1 U104 ( .A(tempResult_adjusted_11_), .B(tempResult_adjusted_12_), .S(
        n8), .Z(result[11]) );
  MUX2_X1 U105 ( .A(tempResult_adjusted_12_), .B(tempResult_adjusted_13_), .S(
        n8), .Z(result[12]) );
  MUX2_X1 U106 ( .A(tempResult_adjusted_13_), .B(tempResult_adjusted_14_), .S(
        n8), .Z(result[13]) );
  MUX2_X1 U107 ( .A(tempResult_adjusted_14_), .B(tempResult_adjusted_15_), .S(
        n8), .Z(result[14]) );
  MUX2_X1 U108 ( .A(tempResult_adjusted_15_), .B(tempResult_adjusted_16_), .S(
        n8), .Z(result[15]) );
  MUX2_X1 U109 ( .A(tempResult_adjusted_16_), .B(tempResult_adjusted_17_), .S(
        n8), .Z(result[16]) );
  MUX2_X1 U110 ( .A(tempResult_adjusted_17_), .B(tempResult_adjusted_18_), .S(
        n8), .Z(result[17]) );
  MUX2_X1 U111 ( .A(tempResult_adjusted_18_), .B(tempResult_adjusted_19_), .S(
        n8), .Z(result[18]) );
  MUX2_X1 U112 ( .A(tempResult_adjusted_19_), .B(tempResult_adjusted_20_), .S(
        n8), .Z(result[19]) );
  MUX2_X1 U113 ( .A(tempResult_adjusted_20_), .B(tempResult_adjusted_21_), .S(
        n8), .Z(result[20]) );
  MUX2_X1 U114 ( .A(tempResult_adjusted_21_), .B(tempResult_adjusted_22_), .S(
        n8), .Z(result[21]) );
  MUX2_X1 U115 ( .A(tempResult_adjusted_22_), .B(tempResult_adjusted_23_), .S(
        n8), .Z(result[22]) );
endmodule


module Normalize ( e, a, cout, normExponent, normResult );
  input [7:0] e;
  input [23:0] a;
  output [7:0] normExponent;
  output [23:0] normResult;
  input cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919;

  OR2_X1 U2 ( .A1(n891), .A2(n706), .ZN(n515) );
  INV_X1 U3 ( .A(n175), .ZN(n906) );
  OR2_X1 U4 ( .A1(n1558), .A2(n441), .ZN(n916) );
  OR2_X1 U5 ( .A1(n218), .A2(n915), .ZN(n774) );
  OR2_X1 U6 ( .A1(n1028), .A2(n263), .ZN(n765) );
  BUF_X1 U7 ( .A(n1204), .Z(n574) );
  AOI211_X1 U8 ( .C1(n1534), .C2(n1248), .A(n646), .B(n1137), .ZN(n1113) );
  AND2_X1 U9 ( .A1(n274), .A2(n1255), .ZN(n677) );
  INV_X1 U10 ( .A(n1567), .ZN(n1681) );
  AOI211_X1 U11 ( .C1(n1540), .C2(n1470), .A(n51), .B(n1337), .ZN(n1313) );
  OAI222_X1 U12 ( .A1(n1705), .A2(n246), .B1(n1722), .B2(n814), .C1(n812), 
        .C2(n1724), .ZN(n1766) );
  INV_X1 U13 ( .A(n1577), .ZN(n1780) );
  OR2_X1 U14 ( .A1(n608), .A2(n375), .ZN(n1488) );
  INV_X1 U15 ( .A(e[6]), .ZN(n727) );
  INV_X1 U16 ( .A(e[1]), .ZN(n302) );
  XNOR2_X1 U17 ( .A(n311), .B(n205), .ZN(n837) );
  OAI222_X1 U18 ( .A1(n1799), .A2(n397), .B1(n1811), .B2(n815), .C1(n823), 
        .C2(n1813), .ZN(n1840) );
  INV_X1 U19 ( .A(n1587), .ZN(n1849) );
  BUF_X2 U20 ( .A(n1870), .Z(n816) );
  OR2_X1 U21 ( .A1(n448), .A2(n1677), .ZN(n1911) );
  INV_X1 U22 ( .A(n728), .ZN(n1) );
  OR2_X1 U23 ( .A1(n2), .A2(n1521), .ZN(n1157) );
  NAND2_X1 U24 ( .A1(n590), .A2(n1), .ZN(n2) );
  AND2_X2 U25 ( .A1(n798), .A2(n528), .ZN(n304) );
  AOI211_X1 U26 ( .C1(n1188), .C2(n1187), .A(n803), .B(n1209), .ZN(n3) );
  OR2_X1 U27 ( .A1(n1543), .A2(n1226), .ZN(n4) );
  NAND2_X1 U28 ( .A1(n4), .A2(n1225), .ZN(n1227) );
  OR2_X1 U29 ( .A1(n224), .A2(n371), .ZN(n5) );
  NAND2_X1 U30 ( .A1(n5), .A2(n669), .ZN(n1127) );
  CLKBUF_X1 U31 ( .A(n621), .Z(n371) );
  OR2_X1 U32 ( .A1(n1069), .A2(n153), .ZN(n342) );
  CLKBUF_X1 U33 ( .A(cout), .Z(n410) );
  CLKBUF_X1 U34 ( .A(n57), .Z(n387) );
  OR2_X2 U35 ( .A1(n853), .A2(n449), .ZN(n833) );
  BUF_X1 U36 ( .A(n983), .Z(n531) );
  OR2_X2 U37 ( .A1(n1454), .A2(n655), .ZN(n1448) );
  OR2_X2 U38 ( .A1(n1523), .A2(n1321), .ZN(n1375) );
  CLKBUF_X1 U39 ( .A(n1720), .Z(n822) );
  XOR2_X1 U40 ( .A(n217), .B(e[7]), .Z(n6) );
  NOR2_X1 U41 ( .A1(n571), .A2(n296), .ZN(n7) );
  CLKBUF_X1 U42 ( .A(n1481), .Z(n30) );
  NOR2_X1 U43 ( .A1(n954), .A2(n951), .ZN(n8) );
  AND2_X1 U44 ( .A1(n247), .A2(n279), .ZN(n9) );
  NOR2_X1 U45 ( .A1(n428), .A2(n765), .ZN(n10) );
  AND2_X1 U46 ( .A1(n1190), .A2(n1207), .ZN(n11) );
  AND2_X1 U47 ( .A1(n1158), .A2(n1162), .ZN(n12) );
  AND2_X1 U48 ( .A1(n1419), .A2(n1401), .ZN(n13) );
  NAND2_X1 U49 ( .A1(n1019), .A2(n1021), .ZN(n14) );
  INV_X1 U50 ( .A(e[2]), .ZN(n205) );
  NOR3_X1 U51 ( .A1(n980), .A2(n990), .A3(n983), .ZN(n229) );
  OAI21_X1 U52 ( .B1(n976), .B2(n182), .A(n17), .ZN(n977) );
  NAND2_X1 U53 ( .A1(n632), .A2(n176), .ZN(n962) );
  NAND4_X1 U54 ( .A1(n9), .A2(n19), .A3(n20), .A4(n18), .ZN(n1037) );
  AOI22_X1 U55 ( .A1(n981), .A2(n188), .B1(n534), .B2(n496), .ZN(n15) );
  INV_X1 U56 ( .A(n15), .ZN(n980) );
  NAND3_X1 U57 ( .A1(n16), .A2(n614), .A3(n690), .ZN(n960) );
  INV_X1 U58 ( .A(n122), .ZN(n16) );
  NAND3_X1 U59 ( .A1(n1042), .A2(n300), .A3(n1043), .ZN(n1038) );
  OAI21_X1 U60 ( .B1(n1027), .B2(n778), .A(n1026), .ZN(n1028) );
  OAI211_X1 U61 ( .C1(n975), .C2(n141), .A(n8), .B(n577), .ZN(n17) );
  INV_X1 U62 ( .A(n17), .ZN(n496) );
  NOR3_X1 U63 ( .A1(n990), .A2(n983), .A3(n980), .ZN(n1007) );
  INV_X1 U64 ( .A(n1028), .ZN(n18) );
  INV_X1 U65 ( .A(n1025), .ZN(n19) );
  INV_X1 U66 ( .A(n1022), .ZN(n20) );
  OAI211_X1 U67 ( .C1(n1254), .C2(n1253), .A(n1312), .B(n809), .ZN(n1553) );
  BUF_X1 U68 ( .A(n1543), .Z(n809) );
  OAI21_X1 U69 ( .B1(n1451), .B2(n58), .A(n671), .ZN(n21) );
  NAND4_X1 U70 ( .A1(n654), .A2(n393), .A3(n1494), .A4(n57), .ZN(n22) );
  AND2_X2 U71 ( .A1(n1898), .A2(n96), .ZN(n94) );
  CLKBUF_X1 U72 ( .A(n666), .Z(n23) );
  INV_X1 U73 ( .A(n1679), .ZN(n666) );
  CLKBUF_X1 U74 ( .A(n1450), .Z(n309) );
  AND2_X1 U75 ( .A1(n1614), .A2(n47), .ZN(n24) );
  OAI21_X1 U76 ( .B1(n1603), .B2(n137), .A(n1602), .ZN(n25) );
  OAI21_X1 U77 ( .B1(n1603), .B2(n137), .A(n1602), .ZN(n1915) );
  INV_X1 U78 ( .A(n1609), .ZN(n26) );
  NOR2_X1 U79 ( .A1(n121), .A2(n1612), .ZN(n27) );
  AND2_X1 U80 ( .A1(n1489), .A2(n28), .ZN(n97) );
  NOR2_X1 U81 ( .A1(n609), .A2(n309), .ZN(n28) );
  OR2_X2 U82 ( .A1(n301), .A2(n148), .ZN(n609) );
  OAI21_X1 U83 ( .B1(n559), .B2(n1593), .A(n1600), .ZN(n29) );
  NAND3_X1 U84 ( .A1(n586), .A2(n1611), .A3(n45), .ZN(n31) );
  NAND3_X1 U85 ( .A1(n1916), .A2(n1915), .A3(n482), .ZN(n32) );
  NAND3_X1 U86 ( .A1(n1916), .A2(n25), .A3(n482), .ZN(n33) );
  CLKBUF_X1 U87 ( .A(n121), .Z(n481) );
  BUF_X1 U88 ( .A(n1598), .Z(n34) );
  XNOR2_X1 U89 ( .A(n587), .B(n103), .ZN(n1916) );
  OR2_X1 U90 ( .A1(n38), .A2(n30), .ZN(n35) );
  OR2_X1 U91 ( .A1(n38), .A2(n30), .ZN(n1596) );
  NOR2_X1 U92 ( .A1(n73), .A2(n650), .ZN(n36) );
  XNOR2_X1 U93 ( .A(n1448), .B(n433), .ZN(n37) );
  OAI21_X1 U94 ( .B1(n31), .B2(n55), .A(n1895), .ZN(n38) );
  OAI21_X1 U95 ( .B1(n1489), .B2(n710), .A(n1488), .ZN(n39) );
  CLKBUF_X1 U96 ( .A(n1478), .Z(n95) );
  CLKBUF_X1 U97 ( .A(n1910), .Z(n40) );
  OAI21_X1 U98 ( .B1(n387), .B2(n1492), .A(n1491), .ZN(n41) );
  AND2_X1 U99 ( .A1(n1486), .A2(n514), .ZN(n45) );
  NAND4_X1 U100 ( .A1(n1484), .A2(n37), .A3(n1480), .A4(n1477), .ZN(n42) );
  OR2_X1 U101 ( .A1(n35), .A2(n95), .ZN(n43) );
  OR2_X1 U102 ( .A1(n49), .A2(n446), .ZN(n44) );
  OAI211_X1 U103 ( .C1(n105), .C2(n101), .A(n1631), .B(n802), .ZN(n46) );
  INV_X1 U104 ( .A(n1490), .ZN(n47) );
  BUF_X1 U105 ( .A(n253), .Z(n48) );
  OR2_X1 U106 ( .A1(n52), .A2(n73), .ZN(n49) );
  OR2_X1 U107 ( .A1(n52), .A2(n73), .ZN(n1479) );
  CLKBUF_X1 U108 ( .A(n1356), .Z(n50) );
  OAI21_X1 U109 ( .B1(n290), .B2(n108), .A(n1350), .ZN(n51) );
  OR2_X1 U110 ( .A1(n313), .A2(n593), .ZN(n201) );
  OR2_X1 U111 ( .A1(n313), .A2(n568), .ZN(n592) );
  OAI211_X1 U112 ( .C1(n1476), .C2(n1475), .A(n1631), .B(n802), .ZN(n52) );
  OAI21_X1 U113 ( .B1(n62), .B2(n1316), .A(n1322), .ZN(n53) );
  OR2_X1 U114 ( .A1(n1668), .A2(n54), .ZN(n1334) );
  OR2_X1 U115 ( .A1(n745), .A2(n233), .ZN(n54) );
  NAND4_X1 U116 ( .A1(n1599), .A2(n1601), .A3(n1594), .A4(n1597), .ZN(n55) );
  CLKBUF_X1 U117 ( .A(n1439), .Z(n148) );
  CLKBUF_X1 U118 ( .A(n1608), .Z(n56) );
  INV_X1 U119 ( .A(n1456), .ZN(n57) );
  INV_X1 U120 ( .A(n417), .ZN(n58) );
  OAI21_X1 U121 ( .B1(n610), .B2(n787), .A(n1293), .ZN(n59) );
  NAND4_X1 U122 ( .A1(n1368), .A2(n244), .A3(n275), .A4(n1362), .ZN(n60) );
  NAND4_X1 U123 ( .A1(n1356), .A2(n1376), .A3(n1371), .A4(n1372), .ZN(n61) );
  CLKBUF_X1 U124 ( .A(n1317), .Z(n62) );
  OAI21_X1 U125 ( .B1(n270), .B2(n32), .A(n1632), .ZN(n63) );
  BUF_X2 U126 ( .A(n110), .Z(n64) );
  INV_X1 U127 ( .A(n1402), .ZN(n65) );
  OAI21_X1 U128 ( .B1(n786), .B2(n1365), .A(n322), .ZN(n66) );
  CLKBUF_X1 U129 ( .A(n1453), .Z(n71) );
  CLKBUF_X1 U130 ( .A(n1401), .Z(n67) );
  INV_X1 U131 ( .A(n447), .ZN(n68) );
  NAND4_X1 U132 ( .A1(n189), .A2(n1335), .A3(n1329), .A4(n78), .ZN(n69) );
  NOR2_X1 U133 ( .A1(n1592), .A2(n104), .ZN(n70) );
  OR2_X1 U134 ( .A1(n1370), .A2(n1369), .ZN(n72) );
  OR2_X1 U135 ( .A1(n1370), .A2(n1369), .ZN(n725) );
  OAI21_X1 U136 ( .B1(n1441), .B2(n801), .A(n1440), .ZN(n73) );
  CLKBUF_X1 U137 ( .A(n1448), .Z(n74) );
  OAI21_X1 U138 ( .B1(n234), .B2(n292), .A(n1325), .ZN(n75) );
  OAI21_X1 U139 ( .B1(n234), .B2(n292), .A(n1325), .ZN(n76) );
  OAI22_X1 U140 ( .A1(n1551), .A2(n139), .B1(n1582), .B2(n268), .ZN(n77) );
  INV_X1 U141 ( .A(n59), .ZN(n78) );
  INV_X1 U142 ( .A(n501), .ZN(n658) );
  XNOR2_X1 U143 ( .A(n546), .B(n613), .ZN(n79) );
  CLKBUF_X1 U144 ( .A(n77), .Z(n80) );
  AND2_X1 U145 ( .A1(n639), .A2(n1285), .ZN(n81) );
  OR2_X1 U146 ( .A1(n242), .A2(n905), .ZN(n82) );
  CLKBUF_X1 U147 ( .A(n698), .Z(n83) );
  NOR2_X1 U148 ( .A1(n699), .A2(n700), .ZN(n698) );
  BUF_X1 U149 ( .A(n1294), .Z(n610) );
  CLKBUF_X1 U150 ( .A(n782), .Z(n84) );
  CLKBUF_X1 U151 ( .A(n1561), .Z(n85) );
  OR2_X1 U152 ( .A1(n82), .A2(n920), .ZN(n86) );
  OAI21_X1 U153 ( .B1(n1362), .B2(n372), .A(n1361), .ZN(n87) );
  AND2_X1 U154 ( .A1(n1614), .A2(n1608), .ZN(n88) );
  NAND2_X1 U155 ( .A1(n673), .A2(n547), .ZN(n89) );
  XOR2_X1 U156 ( .A(n74), .B(n433), .Z(n90) );
  NAND3_X1 U157 ( .A1(n88), .A2(n1611), .A3(n45), .ZN(n91) );
  NAND4_X1 U158 ( .A1(n1317), .A2(n1320), .A3(n1323), .A4(n1324), .ZN(n92) );
  NAND2_X1 U159 ( .A1(n1640), .A2(n93), .ZN(n1444) );
  NOR2_X1 U160 ( .A1(n104), .A2(n1402), .ZN(n93) );
  INV_X1 U161 ( .A(n23), .ZN(n96) );
  NAND2_X1 U162 ( .A1(n36), .A2(n97), .ZN(n1486) );
  AND2_X1 U163 ( .A1(n394), .A2(n714), .ZN(n203) );
  CLKBUF_X1 U164 ( .A(n425), .Z(n98) );
  NOR2_X1 U165 ( .A1(n896), .A2(n893), .ZN(n99) );
  OAI21_X1 U166 ( .B1(n693), .B2(n1418), .A(n1417), .ZN(n100) );
  CLKBUF_X1 U167 ( .A(n1476), .Z(n101) );
  CLKBUF_X1 U168 ( .A(n39), .Z(n102) );
  CLKBUF_X1 U169 ( .A(n1599), .Z(n103) );
  BUF_X1 U170 ( .A(n1405), .Z(n104) );
  NAND4_X1 U171 ( .A1(n1487), .A2(n1489), .A3(n387), .A4(n68), .ZN(n105) );
  CLKBUF_X1 U172 ( .A(n1399), .Z(n368) );
  AOI21_X1 U173 ( .B1(n107), .B2(n490), .A(n693), .ZN(n106) );
  INV_X1 U174 ( .A(n1419), .ZN(n107) );
  OAI21_X1 U175 ( .B1(n290), .B2(n108), .A(n1350), .ZN(n643) );
  NAND4_X1 U176 ( .A1(n287), .A2(n1298), .A3(n1294), .A4(n698), .ZN(n108) );
  NOR2_X1 U177 ( .A1(n1379), .A2(n1378), .ZN(n109) );
  OAI22_X1 U178 ( .A1(n520), .A2(n1678), .B1(n23), .B2(n1896), .ZN(n110) );
  NOR2_X1 U179 ( .A1(n72), .A2(n66), .ZN(n111) );
  OAI21_X1 U180 ( .B1(n1353), .B2(n237), .A(n420), .ZN(n112) );
  OAI21_X1 U181 ( .B1(n264), .B2(n1292), .A(n1291), .ZN(n113) );
  OR2_X1 U182 ( .A1(n1522), .A2(n1259), .ZN(n114) );
  NOR2_X1 U183 ( .A1(n112), .A2(n499), .ZN(n115) );
  AOI211_X1 U184 ( .C1(n466), .C2(n1397), .A(n810), .B(n1420), .ZN(n116) );
  NOR2_X1 U185 ( .A1(n1050), .A2(n536), .ZN(n117) );
  BUF_X1 U186 ( .A(n1049), .Z(n536) );
  OR2_X1 U187 ( .A1(n254), .A2(n132), .ZN(n118) );
  NAND4_X1 U188 ( .A1(n1099), .A2(n1095), .A3(n602), .A4(n1102), .ZN(n119) );
  OAI21_X1 U189 ( .B1(n92), .B2(n1314), .A(n1313), .ZN(n120) );
  OAI21_X1 U190 ( .B1(n607), .B2(n1614), .A(n1613), .ZN(n121) );
  AOI211_X1 U191 ( .C1(n1007), .C2(n1006), .A(n800), .B(n1029), .ZN(n1008) );
  OAI21_X1 U192 ( .B1(n937), .B2(n84), .A(n936), .ZN(n122) );
  OAI21_X1 U193 ( .B1(n1021), .B2(n557), .A(n1020), .ZN(n123) );
  AOI21_X1 U194 ( .B1(n125), .B2(n123), .A(n126), .ZN(n124) );
  NAND2_X1 U195 ( .A1(n308), .A2(n288), .ZN(n125) );
  NOR2_X1 U196 ( .A1(n761), .A2(n191), .ZN(n126) );
  NAND2_X1 U197 ( .A1(n1008), .A2(n286), .ZN(n127) );
  BUF_X1 U198 ( .A(n564), .Z(n755) );
  NAND4_X1 U199 ( .A1(n735), .A2(n240), .A3(n1062), .A4(n1063), .ZN(n128) );
  NAND2_X1 U200 ( .A1(n743), .A2(n129), .ZN(n717) );
  AND2_X1 U201 ( .A1(n1021), .A2(n1019), .ZN(n129) );
  INV_X1 U202 ( .A(n144), .ZN(n130) );
  CLKBUF_X1 U203 ( .A(n1039), .Z(n626) );
  BUF_X1 U204 ( .A(n124), .Z(n754) );
  CLKBUF_X1 U205 ( .A(n239), .Z(n131) );
  OR2_X1 U206 ( .A1(n254), .A2(n132), .ZN(n234) );
  OR2_X1 U207 ( .A1(n255), .A2(n133), .ZN(n132) );
  INV_X1 U208 ( .A(n293), .ZN(n133) );
  OR2_X1 U209 ( .A1(n1026), .A2(n134), .ZN(n279) );
  OR2_X1 U210 ( .A1(n667), .A2(n14), .ZN(n134) );
  NAND2_X1 U211 ( .A1(n552), .A2(n135), .ZN(n756) );
  NOR2_X1 U212 ( .A1(n428), .A2(n757), .ZN(n135) );
  OR2_X1 U213 ( .A1(n891), .A2(n706), .ZN(n136) );
  NAND2_X1 U214 ( .A1(n317), .A2(n455), .ZN(n137) );
  OAI21_X1 U215 ( .B1(n1332), .B2(n543), .A(n347), .ZN(n138) );
  OR4_X1 U216 ( .A1(n962), .A2(n227), .A3(n965), .A4(n967), .ZN(n141) );
  INV_X1 U217 ( .A(n1008), .ZN(n1721) );
  OAI21_X1 U218 ( .B1(n171), .B2(n258), .A(n1313), .ZN(n139) );
  OAI211_X1 U219 ( .C1(n128), .C2(n1057), .A(n805), .B(n1112), .ZN(n140) );
  OR2_X1 U220 ( .A1(n770), .A2(n920), .ZN(n423) );
  OAI21_X2 U221 ( .B1(n953), .B2(n1564), .A(n952), .ZN(n954) );
  OR4_X1 U222 ( .A1(n262), .A2(n912), .A3(n917), .A4(n920), .ZN(n924) );
  INV_X1 U223 ( .A(n153), .ZN(n142) );
  BUF_X1 U224 ( .A(n322), .Z(n143) );
  BUF_X1 U225 ( .A(n944), .Z(n144) );
  CLKBUF_X1 U226 ( .A(n1360), .Z(n316) );
  CLKBUF_X3 U227 ( .A(n1867), .Z(n824) );
  BUF_X1 U228 ( .A(n1331), .Z(n347) );
  XNOR2_X1 U229 ( .A(n145), .B(n292), .ZN(n1371) );
  NOR2_X1 U230 ( .A1(n159), .A2(n254), .ZN(n145) );
  BUF_X1 U231 ( .A(n80), .Z(n730) );
  NOR2_X1 U232 ( .A1(n254), .A2(n255), .ZN(n146) );
  OR2_X1 U233 ( .A1(n1319), .A2(n1286), .ZN(n1322) );
  CLKBUF_X1 U234 ( .A(n644), .Z(n147) );
  NAND2_X1 U235 ( .A1(n222), .A2(n751), .ZN(n1555) );
  CLKBUF_X1 U236 ( .A(n1041), .Z(n162) );
  BUF_X1 U237 ( .A(n1557), .Z(n222) );
  NOR2_X1 U238 ( .A1(n140), .A2(n162), .ZN(n713) );
  BUF_X1 U239 ( .A(n1188), .Z(n476) );
  NAND2_X1 U240 ( .A1(n70), .A2(n500), .ZN(n149) );
  OAI21_X1 U241 ( .B1(n692), .B2(n320), .A(n236), .ZN(n150) );
  OAI21_X1 U242 ( .B1(n924), .B2(n177), .A(n971), .ZN(n151) );
  XNOR2_X1 U243 ( .A(n282), .B(n380), .ZN(n1062) );
  XNOR2_X1 U244 ( .A(n152), .B(n935), .ZN(n956) );
  NOR2_X1 U245 ( .A1(n168), .A2(n773), .ZN(n152) );
  CLKBUF_X1 U246 ( .A(n1047), .Z(n153) );
  INV_X1 U247 ( .A(n340), .ZN(n154) );
  INV_X1 U248 ( .A(n536), .ZN(n155) );
  NOR2_X1 U249 ( .A1(n1557), .A2(n162), .ZN(n411) );
  NOR2_X1 U250 ( .A1(n222), .A2(n156), .ZN(n542) );
  NAND2_X1 U251 ( .A1(n1059), .A2(n755), .ZN(n156) );
  OR2_X1 U252 ( .A1(n665), .A2(n585), .ZN(n157) );
  BUF_X1 U253 ( .A(n1569), .Z(n158) );
  OR2_X1 U254 ( .A1(n255), .A2(n133), .ZN(n159) );
  INV_X1 U255 ( .A(n953), .ZN(n160) );
  OAI21_X1 U256 ( .B1(n929), .B2(n1569), .A(n928), .ZN(n930) );
  OAI21_X1 U257 ( .B1(n744), .B2(n323), .A(n1328), .ZN(n161) );
  BUF_X1 U258 ( .A(n1562), .Z(n199) );
  CLKBUF_X1 U259 ( .A(n911), .Z(n163) );
  BUF_X1 U260 ( .A(n164), .Z(n345) );
  AOI21_X1 U261 ( .B1(n165), .B2(n218), .A(n166), .ZN(n164) );
  NAND2_X1 U262 ( .A1(n766), .A2(n943), .ZN(n165) );
  AND2_X1 U263 ( .A1(n766), .A2(n385), .ZN(n166) );
  NAND2_X1 U264 ( .A1(n738), .A2(n696), .ZN(n167) );
  OR2_X1 U265 ( .A1(n774), .A2(n458), .ZN(n168) );
  NAND3_X1 U266 ( .A1(n907), .A2(n519), .A3(n908), .ZN(n169) );
  OAI21_X1 U267 ( .B1(n1255), .B2(n319), .A(n1260), .ZN(n170) );
  NAND4_X1 U268 ( .A1(n1317), .A2(n1320), .A3(n1323), .A4(n113), .ZN(n171) );
  OAI211_X1 U269 ( .C1(n898), .C2(n899), .A(n946), .B(n804), .ZN(n172) );
  NAND2_X1 U270 ( .A1(n173), .A2(n174), .ZN(n936) );
  NOR2_X1 U271 ( .A1(n86), .A2(n426), .ZN(n173) );
  NOR2_X1 U272 ( .A1(n774), .A2(n458), .ZN(n174) );
  NOR2_X1 U273 ( .A1(n172), .A2(n579), .ZN(n175) );
  OR2_X1 U274 ( .A1(n16), .A2(n202), .ZN(n176) );
  NAND4_X1 U275 ( .A1(n79), .A2(n933), .A3(n926), .A4(n929), .ZN(n177) );
  NAND3_X1 U276 ( .A1(n616), .A2(n914), .A3(n551), .ZN(n178) );
  CLKBUF_X1 U277 ( .A(n964), .Z(n179) );
  OR2_X1 U278 ( .A1(n1562), .A2(n585), .ZN(n180) );
  OR2_X1 U279 ( .A1(n461), .A2(n954), .ZN(n181) );
  NOR2_X1 U280 ( .A1(n1518), .A2(n954), .ZN(n182) );
  OR4_X2 U281 ( .A1(n912), .A2(n262), .A3(n920), .A4(n917), .ZN(n215) );
  OAI21_X1 U282 ( .B1(n280), .B2(n613), .A(n909), .ZN(n183) );
  OAI21_X1 U283 ( .B1(n280), .B2(n613), .A(n909), .ZN(n184) );
  OAI21_X1 U284 ( .B1(n948), .B2(n949), .A(n947), .ZN(n665) );
  AND2_X1 U285 ( .A1(n1021), .A2(n286), .ZN(n185) );
  NAND3_X1 U286 ( .A1(n991), .A2(n532), .A3(n992), .ZN(n186) );
  AND2_X1 U287 ( .A1(n228), .A2(n395), .ZN(n187) );
  OAI21_X1 U288 ( .B1(n203), .B2(n345), .A(n966), .ZN(n188) );
  CLKBUF_X1 U289 ( .A(n1025), .Z(n428) );
  INV_X1 U290 ( .A(n150), .ZN(n189) );
  OR2_X1 U291 ( .A1(n699), .A2(n700), .ZN(n190) );
  AND2_X2 U292 ( .A1(n742), .A2(n1233), .ZN(n633) );
  CLKBUF_X1 U293 ( .A(n762), .Z(n191) );
  OAI21_X1 U294 ( .B1(n996), .B2(n1720), .A(n653), .ZN(n192) );
  OAI21_X1 U295 ( .B1(n215), .B2(n355), .A(n971), .ZN(n193) );
  OAI21_X1 U296 ( .B1(n215), .B2(n355), .A(n971), .ZN(n426) );
  AND2_X1 U297 ( .A1(n225), .A2(n837), .ZN(n194) );
  NOR2_X1 U298 ( .A1(n381), .A2(n503), .ZN(n195) );
  NAND2_X1 U299 ( .A1(n768), .A2(n509), .ZN(n196) );
  INV_X1 U300 ( .A(n157), .ZN(n197) );
  INV_X2 U301 ( .A(n157), .ZN(n198) );
  INV_X1 U302 ( .A(n929), .ZN(n200) );
  OR2_X1 U303 ( .A1(n1091), .A2(n716), .ZN(n707) );
  AND2_X1 U304 ( .A1(n690), .A2(n614), .ZN(n202) );
  BUF_X1 U305 ( .A(n1527), .Z(n813) );
  INV_X1 U306 ( .A(n857), .ZN(n204) );
  NAND2_X1 U307 ( .A1(e[1]), .A2(e[0]), .ZN(n206) );
  NAND2_X1 U308 ( .A1(cout), .A2(n207), .ZN(n310) );
  INV_X1 U309 ( .A(n206), .ZN(n207) );
  BUF_X1 U310 ( .A(n673), .Z(n319) );
  OR2_X1 U311 ( .A1(n833), .A2(n208), .ZN(n847) );
  OR2_X1 U312 ( .A1(n569), .A2(n209), .ZN(n208) );
  INV_X1 U313 ( .A(n216), .ZN(n209) );
  XOR2_X1 U314 ( .A(n1264), .B(n635), .Z(n210) );
  BUF_X1 U315 ( .A(n917), .Z(n218) );
  AND2_X1 U316 ( .A1(n1285), .A2(n221), .ZN(n211) );
  BUF_X1 U317 ( .A(n321), .Z(n212) );
  CLKBUF_X1 U318 ( .A(n287), .Z(n321) );
  NAND2_X1 U319 ( .A1(n394), .A2(n714), .ZN(n213) );
  NAND2_X1 U320 ( .A1(n304), .A2(n573), .ZN(n214) );
  CLKBUF_X1 U321 ( .A(n839), .Z(n216) );
  BUF_X1 U322 ( .A(n776), .Z(n283) );
  AND2_X1 U323 ( .A1(n828), .A2(n421), .ZN(n217) );
  CLKBUF_X1 U324 ( .A(n1297), .Z(n238) );
  NAND4_X1 U325 ( .A1(n567), .A2(n1365), .A3(n1359), .A4(n1362), .ZN(n219) );
  NAND4_X1 U326 ( .A1(n1234), .A2(n1236), .A3(n1238), .A4(n1240), .ZN(n220) );
  AND2_X1 U327 ( .A1(n356), .A2(n269), .ZN(n221) );
  CLKBUF_X1 U328 ( .A(n199), .Z(n223) );
  NOR2_X1 U329 ( .A1(n663), .A2(n369), .ZN(n224) );
  INV_X1 U330 ( .A(n364), .ZN(n225) );
  INV_X1 U331 ( .A(n944), .ZN(n226) );
  OAI21_X1 U332 ( .B1(n203), .B2(n345), .A(n966), .ZN(n227) );
  NOR2_X1 U333 ( .A1(n160), .A2(n665), .ZN(n228) );
  OR2_X1 U334 ( .A1(n1659), .A2(n1089), .ZN(n663) );
  OR2_X1 U335 ( .A1(n364), .A2(n598), .ZN(n230) );
  NOR2_X1 U336 ( .A1(n852), .A2(n851), .ZN(n231) );
  CLKBUF_X1 U337 ( .A(n189), .Z(n543) );
  BUF_X1 U338 ( .A(n1584), .Z(n749) );
  XNOR2_X1 U339 ( .A(n232), .B(n1292), .ZN(n1323) );
  NOR2_X1 U340 ( .A1(n306), .A2(n201), .ZN(n232) );
  OAI21_X1 U341 ( .B1(n81), .B2(n212), .A(n1299), .ZN(n233) );
  INV_X1 U342 ( .A(n1320), .ZN(n235) );
  OR2_X1 U343 ( .A1(n592), .A2(n593), .ZN(n236) );
  NAND4_X1 U344 ( .A1(n1356), .A2(n1376), .A3(n1371), .A4(n1372), .ZN(n237) );
  INV_X1 U345 ( .A(n233), .ZN(n239) );
  INV_X1 U346 ( .A(n1041), .ZN(n240) );
  AND2_X1 U347 ( .A1(n247), .A2(n279), .ZN(n241) );
  OAI21_X1 U348 ( .B1(n900), .B2(n901), .A(n906), .ZN(n242) );
  CLKBUF_X1 U349 ( .A(n834), .Z(n243) );
  INV_X1 U350 ( .A(n1327), .ZN(n244) );
  INV_X1 U351 ( .A(n1721), .ZN(n245) );
  INV_X2 U352 ( .A(n245), .ZN(n246) );
  OR2_X1 U353 ( .A1(n789), .A2(n1019), .ZN(n247) );
  NOR2_X1 U354 ( .A1(n1257), .A2(n589), .ZN(n248) );
  XOR2_X1 U355 ( .A(n342), .B(n659), .Z(n249) );
  CLKBUF_X1 U356 ( .A(n765), .Z(n553) );
  BUF_X4 U357 ( .A(n1723), .Z(n814) );
  AND2_X1 U358 ( .A1(n797), .A2(n1012), .ZN(n250) );
  OR2_X1 U359 ( .A1(n1183), .A2(n1013), .ZN(n251) );
  OR2_X1 U360 ( .A1(n1183), .A2(n1013), .ZN(n761) );
  CLKBUF_X1 U361 ( .A(n1589), .Z(n252) );
  OR2_X1 U362 ( .A1(n651), .A2(n268), .ZN(n253) );
  OR2_X1 U363 ( .A1(n120), .A2(n745), .ZN(n254) );
  NAND2_X1 U364 ( .A1(n323), .A2(n712), .ZN(n255) );
  OR2_X1 U365 ( .A1(n1334), .A2(n256), .ZN(n1328) );
  NAND2_X1 U366 ( .A1(n323), .A2(n543), .ZN(n256) );
  AND2_X1 U367 ( .A1(n623), .A2(n344), .ZN(n602) );
  AND2_X1 U368 ( .A1(n623), .A2(n344), .ZN(n278) );
  OAI21_X1 U369 ( .B1(n974), .B2(n186), .A(n1035), .ZN(n257) );
  NAND4_X1 U370 ( .A1(n1329), .A2(n1335), .A3(n189), .A4(n1326), .ZN(n258) );
  NAND2_X1 U371 ( .A1(e[1]), .A2(e[0]), .ZN(n259) );
  NAND2_X1 U372 ( .A1(cout), .A2(n260), .ZN(n825) );
  INV_X1 U373 ( .A(n259), .ZN(n260) );
  CLKBUF_X1 U374 ( .A(n687), .Z(n261) );
  OAI21_X1 U375 ( .B1(n913), .B2(n400), .A(n545), .ZN(n262) );
  OAI21_X1 U376 ( .B1(n1009), .B2(n784), .A(n1014), .ZN(n263) );
  OR2_X1 U377 ( .A1(n201), .A2(n306), .ZN(n264) );
  OR2_X1 U378 ( .A1(n201), .A2(n306), .ZN(n1293) );
  OR2_X1 U379 ( .A1(n49), .A2(n265), .ZN(n1491) );
  OR2_X1 U380 ( .A1(n446), .A2(n1456), .ZN(n265) );
  NOR2_X1 U381 ( .A1(n269), .A2(n266), .ZN(n779) );
  NAND2_X1 U382 ( .A1(n1255), .A2(n402), .ZN(n266) );
  OR2_X1 U383 ( .A1(n1257), .A2(n589), .ZN(n267) );
  INV_X1 U384 ( .A(n1540), .ZN(n268) );
  INV_X1 U385 ( .A(n274), .ZN(n269) );
  NAND3_X1 U386 ( .A1(n530), .A2(n26), .A3(n1913), .ZN(n270) );
  OR2_X1 U387 ( .A1(n1595), .A2(n34), .ZN(n271) );
  OR2_X1 U388 ( .A1(n359), .A2(n1598), .ZN(n576) );
  BUF_X1 U389 ( .A(n539), .Z(n317) );
  NOR2_X1 U390 ( .A1(n1257), .A2(n589), .ZN(n272) );
  OR2_X1 U391 ( .A1(n699), .A2(n700), .ZN(n273) );
  NOR2_X1 U392 ( .A1(n1553), .A2(n401), .ZN(n274) );
  INV_X1 U393 ( .A(n1333), .ZN(n275) );
  AND2_X1 U394 ( .A1(n283), .A2(n276), .ZN(n744) );
  AND2_X1 U395 ( .A1(n239), .A2(n543), .ZN(n276) );
  OR2_X1 U396 ( .A1(n1522), .A2(n277), .ZN(n1299) );
  NAND2_X1 U397 ( .A1(n211), .A2(n321), .ZN(n277) );
  OR2_X1 U398 ( .A1(n918), .A2(n436), .ZN(n280) );
  AND2_X1 U399 ( .A1(n391), .A2(n1226), .ZN(n281) );
  OR2_X1 U400 ( .A1(n756), .A2(n251), .ZN(n282) );
  OR2_X1 U401 ( .A1(n756), .A2(n761), .ZN(n388) );
  NOR2_X1 U402 ( .A1(n295), .A2(n392), .ZN(n391) );
  CLKBUF_X1 U403 ( .A(n391), .Z(n572) );
  CLKBUF_X1 U404 ( .A(n263), .Z(n284) );
  OAI21_X1 U405 ( .B1(n1009), .B2(n784), .A(n1014), .ZN(n1010) );
  OR2_X1 U406 ( .A1(n1026), .A2(n285), .ZN(n1020) );
  OR2_X1 U407 ( .A1(n535), .A2(n989), .ZN(n285) );
  AND2_X1 U408 ( .A1(n1008), .A2(n286), .ZN(n743) );
  AND2_X1 U409 ( .A1(n307), .A2(n507), .ZN(n286) );
  INV_X1 U410 ( .A(n1270), .ZN(n287) );
  AND2_X1 U411 ( .A1(n1040), .A2(n10), .ZN(n288) );
  NOR2_X1 U412 ( .A1(n289), .A2(n201), .ZN(n787) );
  OR2_X1 U413 ( .A1(n568), .A2(n190), .ZN(n289) );
  OR2_X1 U414 ( .A1(n1011), .A2(n977), .ZN(n1014) );
  NAND3_X1 U415 ( .A1(n210), .A2(n1290), .A3(n588), .ZN(n290) );
  AOI211_X1 U416 ( .C1(n229), .C2(n1006), .A(n800), .B(n1029), .ZN(n291) );
  XNOR2_X1 U417 ( .A(n264), .B(n1292), .ZN(n292) );
  CLKBUF_X1 U418 ( .A(n1326), .Z(n293) );
  AND2_X1 U419 ( .A1(n304), .A2(n574), .ZN(n294) );
  AND2_X1 U420 ( .A1(n1151), .A2(n1191), .ZN(n295) );
  OAI21_X1 U421 ( .B1(n1161), .B2(n1162), .A(n1160), .ZN(n296) );
  NAND2_X1 U422 ( .A1(n672), .A2(n297), .ZN(n1201) );
  AND2_X1 U423 ( .A1(n574), .A2(n1202), .ZN(n297) );
  OR2_X1 U424 ( .A1(n271), .A2(n481), .ZN(n298) );
  NAND2_X1 U425 ( .A1(n291), .A2(n299), .ZN(n1026) );
  AND2_X1 U426 ( .A1(n507), .A2(n1027), .ZN(n299) );
  NOR2_X1 U427 ( .A1(n1010), .A2(n1013), .ZN(n300) );
  NAND2_X1 U428 ( .A1(n1494), .A2(n57), .ZN(n301) );
  XNOR2_X1 U429 ( .A(n303), .B(n302), .ZN(n831) );
  NAND2_X1 U430 ( .A1(n410), .A2(e[0]), .ZN(n303) );
  INV_X1 U431 ( .A(n568), .ZN(n305) );
  NAND2_X1 U432 ( .A1(n597), .A2(n305), .ZN(n306) );
  NOR2_X1 U433 ( .A1(n531), .A2(n535), .ZN(n307) );
  INV_X1 U434 ( .A(n324), .ZN(n308) );
  NAND3_X1 U435 ( .A1(cout), .A2(e[1]), .A3(e[0]), .ZN(n311) );
  OAI211_X1 U436 ( .C1(n105), .C2(n101), .A(n1631), .B(n802), .ZN(n312) );
  OAI21_X1 U437 ( .B1(n1283), .B2(n1284), .A(n1350), .ZN(n313) );
  OAI211_X1 U438 ( .C1(n22), .C2(n42), .A(n1631), .B(n802), .ZN(n650) );
  INV_X1 U439 ( .A(n253), .ZN(n314) );
  INV_X1 U440 ( .A(n48), .ZN(n315) );
  NAND4_X1 U441 ( .A1(n1294), .A2(n287), .A3(n1298), .A4(n698), .ZN(n318) );
  CLKBUF_X1 U442 ( .A(n1154), .Z(n325) );
  CLKBUF_X1 U443 ( .A(n843), .Z(n413) );
  CLKBUF_X1 U444 ( .A(n1298), .Z(n320) );
  OR2_X1 U445 ( .A1(n1364), .A2(n731), .ZN(n322) );
  OR2_X1 U446 ( .A1(n376), .A2(n731), .ZN(n724) );
  AOI222_X1 U447 ( .A1(n730), .A2(n1507), .B1(n315), .B2(n1626), .C1(n1849), 
        .C2(n1394), .ZN(n1395) );
  INV_X1 U448 ( .A(n238), .ZN(n323) );
  OR2_X1 U449 ( .A1(n1403), .A2(n1357), .ZN(n1406) );
  OAI21_X1 U450 ( .B1(n1148), .B2(n1149), .A(n1220), .ZN(n648) );
  OAI21_X1 U451 ( .B1(n1037), .B2(n1038), .A(n1081), .ZN(n324) );
  INV_X1 U452 ( .A(n1095), .ZN(n326) );
  OR2_X1 U453 ( .A1(n1888), .A2(n1798), .ZN(n327) );
  OR2_X1 U454 ( .A1(n1778), .A2(n1886), .ZN(n328) );
  NAND3_X1 U455 ( .A1(n327), .A2(n328), .A3(n1777), .ZN(normResult[10]) );
  CLKBUF_X1 U456 ( .A(n1601), .Z(n329) );
  AND2_X1 U457 ( .A1(n881), .A2(n332), .ZN(n330) );
  NOR2_X1 U458 ( .A1(n331), .A2(n204), .ZN(n485) );
  NAND2_X1 U459 ( .A1(n866), .A2(n509), .ZN(n331) );
  NOR2_X1 U460 ( .A1(n333), .A2(n508), .ZN(n332) );
  NOR2_X1 U461 ( .A1(n857), .A2(n471), .ZN(n333) );
  CLKBUF_X1 U462 ( .A(n231), .Z(n563) );
  OAI21_X1 U463 ( .B1(n866), .B2(n373), .A(n865), .ZN(n334) );
  OAI21_X1 U464 ( .B1(n498), .B2(n783), .A(n487), .ZN(n335) );
  OR2_X1 U465 ( .A1(n1091), .A2(n716), .ZN(n1101) );
  OR2_X1 U466 ( .A1(n887), .A2(n652), .ZN(n336) );
  AND2_X1 U467 ( .A1(n357), .A2(n715), .ZN(n337) );
  NAND3_X1 U468 ( .A1(n249), .A2(n1092), .A3(n537), .ZN(n338) );
  CLKBUF_X1 U469 ( .A(n249), .Z(n339) );
  OAI21_X1 U470 ( .B1(n754), .B2(n733), .A(n612), .ZN(n340) );
  NOR2_X1 U471 ( .A1(n121), .A2(n1612), .ZN(n530) );
  NAND2_X1 U472 ( .A1(n713), .A2(n341), .ZN(n1065) );
  AND2_X1 U473 ( .A1(n656), .A2(n142), .ZN(n341) );
  NOR2_X1 U474 ( .A1(n1050), .A2(n1061), .ZN(n343) );
  OR2_X1 U475 ( .A1(n1061), .A2(n1050), .ZN(n344) );
  OR2_X1 U476 ( .A1(n1659), .A2(n346), .ZN(n1122) );
  OR2_X1 U477 ( .A1(n1089), .A2(n1086), .ZN(n346) );
  NOR2_X1 U478 ( .A1(n310), .A2(n348), .ZN(n794) );
  OR2_X1 U479 ( .A1(n561), .A2(n349), .ZN(n348) );
  INV_X1 U480 ( .A(e[4]), .ZN(n349) );
  CLKBUF_X1 U481 ( .A(n1582), .Z(n350) );
  NOR2_X1 U482 ( .A1(n193), .A2(n351), .ZN(n580) );
  OR2_X1 U483 ( .A1(n423), .A2(n218), .ZN(n351) );
  NOR2_X1 U484 ( .A1(n927), .A2(n930), .ZN(n416) );
  OR2_X1 U485 ( .A1(n1911), .A2(n408), .ZN(n352) );
  OR2_X1 U486 ( .A1(n1911), .A2(n408), .ZN(n1914) );
  OR2_X1 U487 ( .A1(n251), .A2(n756), .ZN(n1046) );
  AND2_X1 U488 ( .A1(n1537), .A2(n353), .ZN(n764) );
  AND2_X1 U489 ( .A1(n1040), .A2(n354), .ZN(n353) );
  INV_X1 U490 ( .A(n553), .ZN(n354) );
  NAND4_X1 U491 ( .A1(n931), .A2(n183), .A3(n926), .A4(n929), .ZN(n355) );
  OR2_X1 U492 ( .A1(n1540), .A2(n1258), .ZN(n356) );
  NAND2_X1 U493 ( .A1(n356), .A2(n269), .ZN(n1259) );
  OR2_X1 U494 ( .A1(n437), .A2(n892), .ZN(n357) );
  CLKBUF_X1 U495 ( .A(n308), .Z(n805) );
  OR2_X1 U496 ( .A1(n592), .A2(n358), .ZN(n1296) );
  OR2_X1 U497 ( .A1(n593), .A2(n273), .ZN(n358) );
  OAI21_X1 U498 ( .B1(n559), .B2(n1593), .A(n1600), .ZN(n359) );
  NOR4_X1 U499 ( .A1(n334), .A2(n335), .A3(n872), .A4(n875), .ZN(n360) );
  NOR4_X1 U500 ( .A1(n868), .A2(n867), .A3(n872), .A4(n875), .ZN(n705) );
  NOR2_X1 U501 ( .A1(n311), .A2(n361), .ZN(n419) );
  OR2_X1 U502 ( .A1(n561), .A2(n452), .ZN(n361) );
  INV_X1 U503 ( .A(n570), .ZN(n362) );
  NOR2_X1 U504 ( .A1(n310), .A2(n205), .ZN(n793) );
  INV_X1 U505 ( .A(n1100), .ZN(n363) );
  OR2_X1 U506 ( .A1(n853), .A2(n449), .ZN(n364) );
  AND2_X1 U507 ( .A1(n180), .A2(n578), .ZN(n365) );
  CLKBUF_X1 U508 ( .A(n1868), .Z(n366) );
  AOI21_X1 U509 ( .B1(n360), .B2(n704), .A(n877), .ZN(n367) );
  INV_X1 U510 ( .A(n368), .ZN(n1868) );
  BUF_X1 U511 ( .A(n508), .Z(n768) );
  OR2_X1 U512 ( .A1(n663), .A2(n369), .ZN(n1128) );
  OR2_X1 U513 ( .A1(n664), .A2(n370), .ZN(n369) );
  INV_X1 U514 ( .A(n363), .ZN(n370) );
  OR2_X1 U515 ( .A1(n1101), .A2(n722), .ZN(n555) );
  OAI222_X1 U516 ( .A1(n1747), .A2(n816), .B1(n824), .B2(n1760), .C1(n1734), 
        .C2(n366), .ZN(n1796) );
  OAI222_X1 U517 ( .A1(n1734), .A2(n816), .B1(n824), .B2(n1747), .C1(n1715), 
        .C2(n366), .ZN(n1776) );
  OR2_X1 U518 ( .A1(n825), .A2(n502), .ZN(n827) );
  NOR2_X1 U519 ( .A1(n422), .A2(n497), .ZN(n372) );
  AND2_X1 U520 ( .A1(n508), .A2(n509), .ZN(n373) );
  NAND2_X1 U521 ( .A1(n740), .A2(n839), .ZN(n374) );
  OR2_X1 U522 ( .A1(n609), .A2(n71), .ZN(n375) );
  NAND2_X1 U523 ( .A1(n115), .A2(n1359), .ZN(n376) );
  BUF_X1 U524 ( .A(n386), .Z(n652) );
  XNOR2_X1 U525 ( .A(n377), .B(n1232), .ZN(n1261) );
  NOR2_X1 U526 ( .A1(n683), .A2(n575), .ZN(n377) );
  INV_X1 U527 ( .A(n749), .ZN(n378) );
  INV_X1 U528 ( .A(n1528), .ZN(n379) );
  CLKBUF_X1 U529 ( .A(n1042), .Z(n380) );
  OAI211_X1 U530 ( .C1(n898), .C2(n169), .A(n946), .B(n804), .ZN(n381) );
  OAI211_X1 U531 ( .C1(n169), .C2(n178), .A(n946), .B(n804), .ZN(n382) );
  OAI211_X1 U532 ( .C1(n899), .C2(n178), .A(n946), .B(n804), .ZN(n1558) );
  NOR2_X1 U533 ( .A1(n1598), .A2(n29), .ZN(n482) );
  BUF_X1 U534 ( .A(n274), .Z(n673) );
  AND2_X1 U535 ( .A1(n468), .A2(n469), .ZN(n383) );
  CLKBUF_X1 U536 ( .A(n1911), .Z(n384) );
  AND2_X1 U537 ( .A1(n943), .A2(n942), .ZN(n385) );
  AND2_X1 U538 ( .A1(n468), .A2(n469), .ZN(n855) );
  INV_X1 U539 ( .A(n602), .ZN(n1074) );
  OAI21_X1 U540 ( .B1(n445), .B2(n889), .A(n888), .ZN(n386) );
  OAI21_X1 U541 ( .B1(n895), .B2(n767), .A(n894), .ZN(n389) );
  NOR2_X1 U542 ( .A1(n257), .A2(n538), .ZN(n390) );
  OR2_X1 U543 ( .A1(n683), .A2(n575), .ZN(n1233) );
  AND2_X1 U544 ( .A1(n522), .A2(n1190), .ZN(n392) );
  INV_X1 U545 ( .A(n1450), .ZN(n393) );
  NOR2_X1 U546 ( .A1(n160), .A2(n1650), .ZN(n394) );
  NAND2_X1 U547 ( .A1(n228), .A2(n395), .ZN(n966) );
  AND2_X1 U548 ( .A1(n345), .A2(n714), .ZN(n395) );
  INV_X1 U549 ( .A(n1810), .ZN(n396) );
  INV_X2 U550 ( .A(n396), .ZN(n397) );
  OR2_X1 U551 ( .A1(n242), .A2(n905), .ZN(n770) );
  CLKBUF_X1 U552 ( .A(n367), .Z(n398) );
  INV_X1 U553 ( .A(n804), .ZN(n399) );
  INV_X1 U554 ( .A(n652), .ZN(n400) );
  INV_X1 U555 ( .A(n1258), .ZN(n401) );
  INV_X1 U556 ( .A(n584), .ZN(n1225) );
  INV_X1 U557 ( .A(n1241), .ZN(n402) );
  AND2_X1 U558 ( .A1(n1103), .A2(n680), .ZN(n403) );
  NOR2_X2 U559 ( .A1(n403), .A2(n1098), .ZN(n624) );
  AND2_X1 U560 ( .A1(n754), .A2(n564), .ZN(n404) );
  NAND2_X1 U561 ( .A1(n691), .A2(n405), .ZN(n685) );
  NOR2_X1 U562 ( .A1(n711), .A2(n1208), .ZN(n405) );
  XNOR2_X1 U563 ( .A(n827), .B(n349), .ZN(n842) );
  OR2_X1 U564 ( .A1(n1888), .A2(n1718), .ZN(n406) );
  OR2_X1 U565 ( .A1(n1704), .A2(n1886), .ZN(n407) );
  NAND3_X1 U566 ( .A1(n406), .A2(n407), .A3(n1703), .ZN(normResult[5]) );
  INV_X1 U567 ( .A(n479), .ZN(n408) );
  NOR2_X1 U568 ( .A1(n149), .A2(n417), .ZN(n409) );
  NAND4_X1 U569 ( .A1(n1102), .A2(n154), .A3(n278), .A4(n1095), .ZN(n412) );
  OAI21_X1 U570 ( .B1(n830), .B2(n829), .A(n876), .ZN(n414) );
  OAI211_X1 U571 ( .C1(n1254), .C2(n1253), .A(n1312), .B(n809), .ZN(n415) );
  BUF_X2 U572 ( .A(n398), .Z(n804) );
  INV_X1 U573 ( .A(n1452), .ZN(n417) );
  INV_X1 U574 ( .A(n846), .ZN(n418) );
  XNOR2_X1 U575 ( .A(n419), .B(e[6]), .ZN(n844) );
  INV_X1 U576 ( .A(n1352), .ZN(n420) );
  AND2_X1 U577 ( .A1(n828), .A2(n421), .ZN(n795) );
  NOR2_X1 U578 ( .A1(n452), .A2(n727), .ZN(n421) );
  BUF_X2 U579 ( .A(n1809), .Z(n823) );
  OAI21_X1 U580 ( .B1(n219), .B2(n61), .A(n420), .ZN(n422) );
  OR2_X1 U581 ( .A1(n426), .A2(n86), .ZN(n773) );
  AOI211_X1 U582 ( .C1(n231), .C2(n855), .A(a[22]), .B(n796), .ZN(n424) );
  OAI21_X1 U583 ( .B1(n924), .B2(n177), .A(n971), .ZN(n425) );
  OR2_X1 U584 ( .A1(n648), .A2(n427), .ZN(n591) );
  OR2_X1 U585 ( .A1(n728), .A2(n1136), .ZN(n427) );
  OAI21_X1 U586 ( .B1(n215), .B2(n925), .A(n971), .ZN(n1517) );
  BUF_X1 U587 ( .A(n250), .Z(n784) );
  OR2_X1 U588 ( .A1(n556), .A2(n429), .ZN(n448) );
  NAND2_X1 U589 ( .A1(n26), .A2(n1907), .ZN(n429) );
  NAND2_X1 U590 ( .A1(n317), .A2(n430), .ZN(n1604) );
  AND2_X1 U591 ( .A1(n480), .A2(n431), .ZN(n430) );
  INV_X1 U592 ( .A(n595), .ZN(n431) );
  NAND4_X1 U593 ( .A1(n1443), .A2(n1441), .A3(n1438), .A4(n1445), .ZN(n432) );
  CLKBUF_X1 U594 ( .A(n1443), .Z(n433) );
  NAND2_X1 U595 ( .A1(n357), .A2(n715), .ZN(n434) );
  OR2_X1 U596 ( .A1(n437), .A2(n892), .ZN(n435) );
  NAND2_X1 U597 ( .A1(n435), .A2(n715), .ZN(n893) );
  OR2_X1 U598 ( .A1(n918), .A2(n436), .ZN(n910) );
  OR2_X1 U599 ( .A1(n434), .A2(n336), .ZN(n436) );
  AND2_X1 U600 ( .A1(n703), .A2(n523), .ZN(n437) );
  AND2_X1 U601 ( .A1(n703), .A2(n523), .ZN(n734) );
  NAND3_X1 U602 ( .A1(n416), .A2(n956), .A3(n957), .ZN(n949) );
  INV_X1 U603 ( .A(n585), .ZN(n438) );
  OR2_X1 U604 ( .A1(n381), .A2(n439), .ZN(n545) );
  OR2_X1 U605 ( .A1(n441), .A2(n652), .ZN(n439) );
  OR2_X1 U606 ( .A1(n382), .A2(n503), .ZN(n440) );
  OR2_X1 U607 ( .A1(n579), .A2(n747), .ZN(n441) );
  NOR2_X1 U608 ( .A1(n1650), .A2(n160), .ZN(n690) );
  BUF_X4 U609 ( .A(n1812), .Z(n815) );
  OR2_X1 U610 ( .A1(n858), .A2(n450), .ZN(n873) );
  AND2_X1 U611 ( .A1(n474), .A2(n806), .ZN(n442) );
  OR2_X1 U612 ( .A1(n1888), .A2(n1763), .ZN(n443) );
  OR2_X1 U613 ( .A1(n1750), .A2(n1886), .ZN(n444) );
  NAND3_X1 U614 ( .A1(n443), .A2(n444), .A3(n1749), .ZN(normResult[8]) );
  BUF_X1 U615 ( .A(n63), .Z(n520) );
  AND2_X1 U616 ( .A1(n734), .A2(n892), .ZN(n445) );
  OR2_X1 U617 ( .A1(n1479), .A2(n446), .ZN(n1493) );
  OR2_X1 U618 ( .A1(n148), .A2(n447), .ZN(n446) );
  INV_X1 U619 ( .A(n1494), .ZN(n447) );
  OR2_X1 U620 ( .A1(n832), .A2(n850), .ZN(n851) );
  NAND2_X1 U621 ( .A1(n849), .A2(n831), .ZN(n449) );
  OR2_X1 U622 ( .A1(n204), .A2(n838), .ZN(n450) );
  NAND2_X1 U623 ( .A1(n703), .A2(n451), .ZN(n891) );
  AND2_X1 U624 ( .A1(n523), .A2(n892), .ZN(n451) );
  OAI222_X1 U625 ( .A1(n1871), .A2(n816), .B1(n1869), .B2(n366), .C1(n824), 
        .C2(n1866), .ZN(n1893) );
  INV_X1 U626 ( .A(n1528), .ZN(n585) );
  NAND2_X1 U627 ( .A1(e[4]), .A2(e[5]), .ZN(n452) );
  CLKBUF_X1 U628 ( .A(n1015), .Z(n453) );
  INV_X1 U629 ( .A(n480), .ZN(n454) );
  NAND2_X1 U630 ( .A1(n317), .A2(n455), .ZN(n587) );
  NOR2_X1 U631 ( .A1(n595), .A2(n454), .ZN(n455) );
  INV_X1 U632 ( .A(n609), .ZN(n456) );
  NOR2_X1 U633 ( .A1(n457), .A2(n49), .ZN(n777) );
  NAND2_X1 U634 ( .A1(n1489), .A2(n456), .ZN(n457) );
  INV_X1 U635 ( .A(n937), .ZN(n458) );
  NAND2_X1 U636 ( .A1(n459), .A2(n460), .ZN(n538) );
  NOR2_X1 U637 ( .A1(n954), .A2(n188), .ZN(n459) );
  NOR2_X1 U638 ( .A1(n951), .A2(n533), .ZN(n460) );
  OR2_X1 U639 ( .A1(n181), .A2(n799), .ZN(n981) );
  OR2_X1 U640 ( .A1(n951), .A2(n533), .ZN(n461) );
  INV_X1 U641 ( .A(n442), .ZN(n462) );
  OR2_X1 U642 ( .A1(n1888), .A2(n1750), .ZN(n463) );
  OR2_X1 U643 ( .A1(n1737), .A2(n1886), .ZN(n464) );
  NAND3_X1 U644 ( .A1(n463), .A2(n464), .A3(n1736), .ZN(normResult[7]) );
  NAND2_X2 U645 ( .A1(n96), .A2(n478), .ZN(n1886) );
  NOR2_X1 U646 ( .A1(n495), .A2(n843), .ZN(n465) );
  CLKBUF_X1 U647 ( .A(n1200), .Z(n575) );
  NOR2_X1 U648 ( .A1(n548), .A2(n725), .ZN(n466) );
  NAND4_X1 U649 ( .A1(n1455), .A2(n1452), .A3(n1449), .A4(n489), .ZN(n467) );
  OR2_X1 U650 ( .A1(n1399), .A2(n810), .ZN(n1870) );
  NOR2_X1 U651 ( .A1(n835), .A2(n838), .ZN(n468) );
  NOR2_X1 U652 ( .A1(n840), .A2(n843), .ZN(n469) );
  OAI21_X1 U653 ( .B1(n974), .B2(n186), .A(n1035), .ZN(n470) );
  AND2_X1 U654 ( .A1(n424), .A2(n859), .ZN(n471) );
  OAI21_X1 U655 ( .B1(n294), .B2(n1202), .A(n1201), .ZN(n472) );
  NAND4_X1 U656 ( .A1(n363), .A2(n621), .A3(n624), .A4(n1135), .ZN(n473) );
  OAI21_X1 U657 ( .B1(n33), .B2(n1633), .A(n1632), .ZN(n474) );
  CLKBUF_X1 U658 ( .A(n1582), .Z(n475) );
  OAI21_X1 U659 ( .B1(n467), .B2(n432), .A(n1512), .ZN(n477) );
  OAI21_X1 U660 ( .B1(n91), .B2(n55), .A(n1895), .ZN(n478) );
  OAI21_X1 U661 ( .B1(n270), .B2(n1634), .A(n1632), .ZN(n1677) );
  OAI21_X1 U662 ( .B1(n1514), .B2(n1515), .A(n1895), .ZN(n1672) );
  CLKBUF_X1 U663 ( .A(n1913), .Z(n479) );
  CLKBUF_X1 U664 ( .A(n1611), .Z(n480) );
  INV_X1 U665 ( .A(n889), .ZN(n483) );
  OAI21_X1 U666 ( .B1(n498), .B2(n783), .A(n196), .ZN(n868) );
  OAI21_X1 U667 ( .B1(n881), .B2(n804), .A(n880), .ZN(n484) );
  NAND2_X1 U668 ( .A1(n884), .A2(n330), .ZN(n518) );
  CLKBUF_X1 U669 ( .A(n861), .Z(n486) );
  NAND2_X1 U670 ( .A1(n768), .A2(n509), .ZN(n487) );
  AND2_X1 U671 ( .A1(n808), .A2(n506), .ZN(n637) );
  AOI211_X1 U672 ( .C1(n1398), .C2(n109), .A(n810), .B(n1420), .ZN(n1399) );
  CLKBUF_X1 U673 ( .A(n1455), .Z(n488) );
  AOI21_X1 U674 ( .B1(n107), .B2(n490), .A(n693), .ZN(n489) );
  NAND2_X1 U675 ( .A1(n1400), .A2(n67), .ZN(n490) );
  AND2_X1 U676 ( .A1(n116), .A2(n491), .ZN(n617) );
  AND2_X1 U677 ( .A1(n506), .A2(n1418), .ZN(n491) );
  AND2_X1 U678 ( .A1(n637), .A2(n1418), .ZN(n492) );
  OAI21_X1 U679 ( .B1(n1365), .B2(n786), .A(n143), .ZN(n493) );
  CLKBUF_X1 U680 ( .A(n1512), .Z(n494) );
  OAI21_X1 U681 ( .B1(n243), .B2(n194), .A(n230), .ZN(n495) );
  XNOR2_X1 U682 ( .A(n847), .B(n418), .ZN(n861) );
  OR2_X1 U683 ( .A1(n422), .A2(n497), .ZN(n1358) );
  OR2_X1 U684 ( .A1(n1321), .A2(n53), .ZN(n497) );
  NOR2_X1 U685 ( .A1(n873), .A2(n527), .ZN(n498) );
  OR2_X1 U686 ( .A1(n662), .A2(n1321), .ZN(n499) );
  AND2_X1 U687 ( .A1(n488), .A2(n505), .ZN(n500) );
  NAND2_X1 U688 ( .A1(n70), .A2(n505), .ZN(n501) );
  OAI21_X1 U689 ( .B1(n195), .B2(n337), .A(n916), .ZN(n917) );
  AOI21_X1 U690 ( .B1(n705), .B2(n704), .A(n877), .ZN(n703) );
  NAND2_X1 U691 ( .A1(e[2]), .A2(e[3]), .ZN(n502) );
  OR2_X1 U692 ( .A1(n1558), .A2(n503), .ZN(n918) );
  OR2_X1 U693 ( .A1(n579), .A2(n389), .ZN(n503) );
  NOR2_X1 U694 ( .A1(n1592), .A2(n104), .ZN(n504) );
  AND2_X1 U695 ( .A1(n106), .A2(n65), .ZN(n505) );
  AND2_X1 U696 ( .A1(n1404), .A2(n13), .ZN(n506) );
  AND2_X1 U697 ( .A1(n291), .A2(n507), .ZN(n778) );
  AND2_X1 U698 ( .A1(n1012), .A2(n1009), .ZN(n507) );
  NOR2_X1 U699 ( .A1(n858), .A2(n204), .ZN(n508) );
  AND2_X1 U700 ( .A1(n465), .A2(n874), .ZN(n509) );
  INV_X1 U701 ( .A(n1157), .ZN(n510) );
  AND2_X1 U702 ( .A1(n1161), .A2(n1162), .ZN(n511) );
  INV_X1 U703 ( .A(n1221), .ZN(n512) );
  NAND2_X1 U704 ( .A1(n544), .A2(n590), .ZN(n513) );
  OR2_X1 U705 ( .A1(n1154), .A2(n1156), .ZN(n1164) );
  OR2_X1 U706 ( .A1(n777), .A2(n1487), .ZN(n514) );
  XNOR2_X1 U707 ( .A(n1448), .B(n433), .ZN(n1483) );
  NOR2_X1 U708 ( .A1(n483), .A2(n891), .ZN(n516) );
  OR2_X1 U709 ( .A1(n891), .A2(n483), .ZN(n888) );
  NOR2_X1 U710 ( .A1(n879), .A2(n882), .ZN(n519) );
  NOR2_X1 U711 ( .A1(n518), .A2(n517), .ZN(n704) );
  AND2_X1 U712 ( .A1(n719), .A2(n720), .ZN(n517) );
  OR2_X1 U713 ( .A1(n1610), .A2(n102), .ZN(n1606) );
  NOR2_X1 U714 ( .A1(n825), .A2(n561), .ZN(n828) );
  AND2_X1 U715 ( .A1(n615), .A2(n1418), .ZN(n521) );
  AND2_X1 U716 ( .A1(n798), .A2(n1192), .ZN(n522) );
  AND2_X1 U717 ( .A1(n526), .A2(n895), .ZN(n523) );
  AOI211_X1 U718 ( .C1(n476), .C2(n723), .A(n803), .B(n1209), .ZN(n1189) );
  AND2_X1 U719 ( .A1(n1526), .A2(n849), .ZN(n524) );
  AND2_X1 U720 ( .A1(n639), .A2(n1285), .ZN(n525) );
  NAND2_X1 U721 ( .A1(n367), .A2(n526), .ZN(n883) );
  AND2_X1 U722 ( .A1(n881), .A2(n332), .ZN(n526) );
  INV_X1 U723 ( .A(n871), .ZN(n527) );
  AND2_X1 U724 ( .A1(n3), .A2(n528), .ZN(n672) );
  AND2_X1 U725 ( .A1(n1192), .A2(n11), .ZN(n528) );
  OAI21_X1 U726 ( .B1(n739), .B2(n243), .A(n230), .ZN(n835) );
  OAI21_X1 U727 ( .B1(n1114), .B2(n1115), .A(n1113), .ZN(n529) );
  AOI211_X1 U728 ( .C1(n563), .C2(n855), .A(a[22]), .B(n796), .ZN(n856) );
  BUF_X1 U729 ( .A(n1641), .Z(n806) );
  NOR2_X1 U730 ( .A1(n951), .A2(n954), .ZN(n532) );
  OAI21_X1 U731 ( .B1(n611), .B2(n130), .A(n213), .ZN(n533) );
  NAND2_X1 U732 ( .A1(n496), .A2(n534), .ZN(n984) );
  NOR2_X1 U733 ( .A1(n188), .A2(n533), .ZN(n534) );
  OAI21_X1 U734 ( .B1(n979), .B2(n978), .A(n984), .ZN(n535) );
  NOR2_X1 U735 ( .A1(n1060), .A2(n1058), .ZN(n537) );
  NOR2_X1 U736 ( .A1(n1672), .A2(n540), .ZN(n539) );
  OR2_X1 U737 ( .A1(n560), .A2(n30), .ZN(n540) );
  INV_X1 U738 ( .A(n1564), .ZN(n541) );
  NOR2_X1 U739 ( .A1(n470), .A2(n538), .ZN(n738) );
  NAND2_X1 U740 ( .A1(n544), .A2(n590), .ZN(n1169) );
  AND2_X1 U741 ( .A1(n726), .A2(n12), .ZN(n544) );
  XNOR2_X1 U742 ( .A(n546), .B(n613), .ZN(n931) );
  NOR2_X1 U743 ( .A1(n918), .A2(n606), .ZN(n546) );
  OR2_X1 U744 ( .A1(n382), .A2(n484), .ZN(n903) );
  XNOR2_X1 U745 ( .A(n1411), .B(n550), .ZN(n1443) );
  NAND2_X1 U746 ( .A1(n673), .A2(n547), .ZN(n1264) );
  NOR2_X1 U747 ( .A1(n589), .A2(n769), .ZN(n547) );
  OR2_X1 U748 ( .A1(n1553), .A2(n401), .ZN(n1257) );
  OAI21_X1 U749 ( .B1(n786), .B2(n1365), .A(n322), .ZN(n548) );
  OAI21_X1 U750 ( .B1(n1374), .B2(n143), .A(n1373), .ZN(n549) );
  CLKBUF_X1 U751 ( .A(n1407), .Z(n550) );
  NOR2_X1 U752 ( .A1(n896), .A2(n893), .ZN(n551) );
  OR2_X1 U753 ( .A1(n977), .A2(n997), .ZN(n998) );
  XNOR2_X1 U754 ( .A(n995), .B(n638), .ZN(n1015) );
  NAND2_X1 U755 ( .A1(n552), .A2(n19), .ZN(n762) );
  NOR2_X1 U756 ( .A1(n765), .A2(n123), .ZN(n552) );
  OR2_X1 U757 ( .A1(n1520), .A2(n599), .ZN(n554) );
  OR2_X1 U758 ( .A1(n1520), .A2(n599), .ZN(n1091) );
  OR2_X1 U759 ( .A1(n474), .A2(n34), .ZN(n1900) );
  OR2_X1 U760 ( .A1(n474), .A2(n271), .ZN(n1903) );
  NOR2_X1 U761 ( .A1(n474), .A2(n298), .ZN(n594) );
  OR2_X1 U762 ( .A1(n576), .A2(n121), .ZN(n556) );
  NOR2_X1 U763 ( .A1(n1026), .A2(n667), .ZN(n557) );
  CLKBUF_X1 U764 ( .A(n1574), .Z(n558) );
  NAND3_X1 U765 ( .A1(n1913), .A2(n1910), .A3(n27), .ZN(n1633) );
  INV_X1 U766 ( .A(n95), .ZN(n559) );
  OR2_X1 U767 ( .A1(n35), .A2(n560), .ZN(n1613) );
  NAND2_X1 U768 ( .A1(n1594), .A2(n1614), .ZN(n560) );
  NAND2_X1 U769 ( .A1(e[2]), .A2(e[3]), .ZN(n561) );
  OAI21_X1 U770 ( .B1(n985), .B2(n697), .A(n167), .ZN(n562) );
  AOI21_X1 U771 ( .B1(n284), .B2(n626), .A(n736), .ZN(n564) );
  NOR2_X1 U772 ( .A1(n662), .A2(n1375), .ZN(n565) );
  NAND2_X1 U773 ( .A1(n565), .A2(n566), .ZN(n1366) );
  AND2_X1 U774 ( .A1(n567), .A2(n275), .ZN(n566) );
  INV_X1 U775 ( .A(n161), .ZN(n567) );
  NAND3_X1 U776 ( .A1(n911), .A2(n914), .A3(n99), .ZN(n898) );
  NAND2_X1 U777 ( .A1(n1285), .A2(n221), .ZN(n568) );
  NOR2_X1 U778 ( .A1(n833), .A2(n569), .ZN(n740) );
  OR2_X1 U779 ( .A1(n570), .A2(n598), .ZN(n569) );
  INV_X1 U780 ( .A(n842), .ZN(n570) );
  OAI21_X1 U781 ( .B1(n1158), .B2(n511), .A(n513), .ZN(n571) );
  NAND2_X1 U782 ( .A1(n304), .A2(n573), .ZN(n1198) );
  AND2_X1 U783 ( .A1(n574), .A2(n7), .ZN(n573) );
  NAND3_X1 U784 ( .A1(n1228), .A2(n1230), .A3(n281), .ZN(n1223) );
  INV_X1 U785 ( .A(n973), .ZN(n577) );
  OR2_X1 U786 ( .A1(n1650), .A2(n85), .ZN(n578) );
  NAND2_X1 U787 ( .A1(n180), .A2(n578), .ZN(n1683) );
  OR2_X1 U788 ( .A1(n879), .A2(n882), .ZN(n579) );
  CLKBUF_X1 U789 ( .A(n1236), .Z(n581) );
  CLKBUF_X1 U790 ( .A(n420), .Z(n582) );
  AND2_X1 U791 ( .A1(n708), .A2(n583), .ZN(n684) );
  AND2_X1 U792 ( .A1(n1240), .A2(n1238), .ZN(n583) );
  CLKBUF_X1 U793 ( .A(n261), .Z(n686) );
  NOR2_X1 U794 ( .A1(n681), .A2(n1193), .ZN(n584) );
  AND2_X1 U795 ( .A1(n1614), .A2(n47), .ZN(n586) );
  OR2_X1 U796 ( .A1(n1360), .A2(n1363), .ZN(n1370) );
  NOR2_X1 U797 ( .A1(n1610), .A2(n102), .ZN(n709) );
  NOR2_X1 U798 ( .A1(n1256), .A2(n1259), .ZN(n588) );
  NAND2_X1 U799 ( .A1(n1255), .A2(n603), .ZN(n589) );
  INV_X1 U800 ( .A(n591), .ZN(n601) );
  AND2_X1 U801 ( .A1(n1153), .A2(n1155), .ZN(n590) );
  OR2_X1 U802 ( .A1(n1267), .A2(n1270), .ZN(n593) );
  NAND2_X1 U803 ( .A1(n1608), .A2(n45), .ZN(n595) );
  NOR2_X1 U804 ( .A1(n593), .A2(n592), .ZN(n596) );
  AND2_X1 U805 ( .A1(n610), .A2(n83), .ZN(n597) );
  NOR2_X1 U806 ( .A1(n833), .A2(n598), .ZN(n618) );
  NAND2_X1 U807 ( .A1(n834), .A2(n837), .ZN(n598) );
  OR2_X1 U808 ( .A1(n1060), .A2(n1058), .ZN(n599) );
  OR2_X1 U809 ( .A1(n726), .A2(n1155), .ZN(n600) );
  NAND2_X1 U810 ( .A1(n591), .A2(n600), .ZN(n1156) );
  INV_X1 U811 ( .A(n492), .ZN(n1417) );
  AOI222_X1 U812 ( .A1(n695), .A2(n1076), .B1(n198), .B2(n1107), .C1(n1681), 
        .C2(n1003), .ZN(n1004) );
  INV_X1 U813 ( .A(n394), .ZN(n952) );
  XOR2_X1 U814 ( .A(n1914), .B(n647), .Z(normExponent[6]) );
  AND2_X1 U815 ( .A1(n261), .A2(n402), .ZN(n603) );
  NAND3_X1 U816 ( .A1(n24), .A2(n1611), .A3(n45), .ZN(n1514) );
  INV_X1 U817 ( .A(n664), .ZN(n604) );
  NOR2_X1 U818 ( .A1(n605), .A2(n663), .ZN(n668) );
  NAND2_X1 U819 ( .A1(n670), .A2(n604), .ZN(n605) );
  OR2_X1 U820 ( .A1(n434), .A2(n336), .ZN(n606) );
  NOR2_X1 U821 ( .A1(n95), .A2(n35), .ZN(n607) );
  OR2_X1 U822 ( .A1(n650), .A2(n73), .ZN(n608) );
  NOR2_X1 U823 ( .A1(n608), .A2(n609), .ZN(n710) );
  AND2_X1 U824 ( .A1(n690), .A2(n950), .ZN(n611) );
  INV_X1 U825 ( .A(n1066), .ZN(n612) );
  NAND3_X1 U826 ( .A1(n907), .A2(n519), .A3(n908), .ZN(n899) );
  XNOR2_X1 U827 ( .A(n515), .B(n675), .ZN(n613) );
  NAND2_X1 U828 ( .A1(n690), .A2(n614), .ZN(n963) );
  AND2_X1 U829 ( .A1(n714), .A2(n741), .ZN(n614) );
  AND2_X1 U830 ( .A1(n1412), .A2(n1415), .ZN(n615) );
  INV_X1 U831 ( .A(n887), .ZN(n616) );
  INV_X1 U832 ( .A(n636), .ZN(n1440) );
  OR2_X1 U833 ( .A1(n1393), .A2(n685), .ZN(n683) );
  CLKBUF_X1 U834 ( .A(n1572), .Z(n619) );
  INV_X1 U835 ( .A(n558), .ZN(n620) );
  INV_X1 U836 ( .A(n1096), .ZN(n621) );
  BUF_X1 U837 ( .A(n1105), .Z(n622) );
  OR2_X1 U838 ( .A1(n542), .A2(n752), .ZN(n623) );
  NOR2_X1 U839 ( .A1(n1119), .A2(n664), .ZN(n625) );
  OR2_X1 U840 ( .A1(n1101), .A2(n627), .ZN(n660) );
  OR2_X1 U841 ( .A1(n628), .A2(n326), .ZN(n627) );
  INV_X1 U842 ( .A(n154), .ZN(n628) );
  CLKBUF_X1 U843 ( .A(n1123), .Z(n629) );
  AOI21_X1 U844 ( .B1(n753), .B2(n1028), .A(n759), .ZN(n630) );
  OAI21_X1 U845 ( .B1(n733), .B2(n754), .A(n612), .ZN(n1070) );
  OAI22_X1 U846 ( .A1(n1555), .A2(n620), .B1(n147), .B2(n1572), .ZN(n631) );
  OR2_X1 U847 ( .A1(n963), .A2(n122), .ZN(n632) );
  OR2_X1 U848 ( .A1(n683), .A2(n575), .ZN(n634) );
  XNOR2_X1 U849 ( .A(n634), .B(n1232), .ZN(n635) );
  NOR2_X1 U850 ( .A1(n104), .A2(n477), .ZN(n636) );
  CLKBUF_X1 U851 ( .A(n991), .Z(n638) );
  NOR2_X1 U852 ( .A1(n1522), .A2(n1259), .ZN(n639) );
  NOR2_X1 U853 ( .A1(n1203), .A2(n296), .ZN(n676) );
  NOR2_X1 U854 ( .A1(n1523), .A2(n499), .ZN(n657) );
  AND2_X1 U855 ( .A1(n1574), .A2(n1534), .ZN(n792) );
  INV_X1 U856 ( .A(n792), .ZN(n640) );
  INV_X2 U857 ( .A(n640), .ZN(n641) );
  INV_X1 U858 ( .A(n657), .ZN(n1361) );
  INV_X1 U859 ( .A(n304), .ZN(n1206) );
  INV_X1 U860 ( .A(n801), .ZN(n642) );
  NAND3_X1 U861 ( .A1(n991), .A2(n992), .A3(n532), .ZN(n975) );
  INV_X1 U862 ( .A(n1534), .ZN(n644) );
  OAI21_X1 U863 ( .B1(n412), .B2(n338), .A(n1145), .ZN(n645) );
  OAI21_X1 U864 ( .B1(n338), .B2(n119), .A(n1145), .ZN(n646) );
  CLKBUF_X1 U865 ( .A(n1916), .Z(n647) );
  CLKBUF_X1 U866 ( .A(n956), .Z(n649) );
  BUF_X2 U867 ( .A(n1640), .Z(n801) );
  OAI21_X1 U868 ( .B1(n318), .B2(n1284), .A(n1350), .ZN(n1522) );
  OAI211_X1 U869 ( .C1(n128), .C2(n1057), .A(n805), .B(n1112), .ZN(n1557) );
  OAI21_X1 U870 ( .B1(n1084), .B2(n1083), .A(n1145), .ZN(n1520) );
  OAI21_X1 U871 ( .B1(n171), .B2(n258), .A(n1313), .ZN(n651) );
  OAI21_X1 U872 ( .B1(n1315), .B2(n69), .A(n1313), .ZN(n1668) );
  XNOR2_X1 U873 ( .A(n660), .B(n339), .ZN(n1123) );
  OR2_X1 U874 ( .A1(n707), .A2(n628), .ZN(n1097) );
  INV_X1 U875 ( .A(n182), .ZN(n653) );
  OR2_X1 U876 ( .A1(n986), .A2(n989), .ZN(n990) );
  INV_X1 U877 ( .A(n21), .ZN(n654) );
  OR2_X1 U878 ( .A1(n1416), .A2(n1413), .ZN(n655) );
  NAND2_X1 U879 ( .A1(n411), .A2(n656), .ZN(n1069) );
  AND2_X1 U880 ( .A1(n781), .A2(n404), .ZN(n656) );
  NAND3_X1 U881 ( .A1(n1090), .A2(n1092), .A3(n537), .ZN(n1084) );
  XNOR2_X1 U882 ( .A(n1046), .B(n1045), .ZN(n659) );
  XNOR2_X1 U883 ( .A(n717), .B(n453), .ZN(n1042) );
  NOR2_X1 U884 ( .A1(n1122), .A2(n622), .ZN(n661) );
  OR2_X1 U885 ( .A1(n1318), .A2(n1336), .ZN(n662) );
  OR2_X1 U886 ( .A1(n1122), .A2(n622), .ZN(n1133) );
  OR2_X1 U887 ( .A1(n701), .A2(n1086), .ZN(n664) );
  NAND2_X1 U888 ( .A1(n308), .A2(n288), .ZN(n1048) );
  OR2_X1 U889 ( .A1(n1596), .A2(n95), .ZN(n1600) );
  INV_X1 U890 ( .A(n1024), .ZN(n667) );
  OAI21_X1 U891 ( .B1(n948), .B2(n949), .A(n947), .ZN(n1650) );
  XNOR2_X1 U892 ( .A(n668), .B(n1126), .ZN(n1165) );
  OR4_X2 U893 ( .A1(n1127), .A2(n1132), .A3(n1130), .A4(n1136), .ZN(n1148) );
  AOI222_X1 U894 ( .A1(n679), .A2(n1277), .B1(n641), .B2(n1307), .C1(n1780), 
        .C2(n1184), .ZN(n1185) );
  NAND2_X1 U895 ( .A1(n625), .A2(n670), .ZN(n669) );
  AND2_X1 U896 ( .A1(n371), .A2(n363), .ZN(n670) );
  OR2_X1 U897 ( .A1(n1454), .A2(n655), .ZN(n674) );
  OR2_X1 U898 ( .A1(n1454), .A2(n417), .ZN(n671) );
  AND2_X1 U899 ( .A1(n719), .A2(n720), .ZN(n675) );
  INV_X1 U900 ( .A(n677), .ZN(n1260) );
  INV_X1 U901 ( .A(n625), .ZN(n1131) );
  OAI21_X1 U902 ( .B1(n473), .B2(n1115), .A(n1113), .ZN(n1659) );
  INV_X1 U903 ( .A(n631), .ZN(n678) );
  INV_X1 U904 ( .A(n678), .ZN(n679) );
  XNOR2_X1 U905 ( .A(n1169), .B(n1165), .ZN(n1194) );
  INV_X1 U906 ( .A(n1102), .ZN(n680) );
  NAND2_X1 U907 ( .A1(n1235), .A2(n575), .ZN(n742) );
  OAI21_X1 U908 ( .B1(n220), .B2(n1223), .A(n512), .ZN(n681) );
  INV_X1 U909 ( .A(n809), .ZN(n682) );
  OAI21_X1 U910 ( .B1(n1222), .B2(n1223), .A(n512), .ZN(n1393) );
  OR2_X1 U911 ( .A1(n681), .A2(n685), .ZN(n1235) );
  AOI21_X1 U912 ( .B1(n1239), .B2(n1205), .A(n684), .ZN(n687) );
  NOR2_X1 U913 ( .A1(n1224), .A2(n1227), .ZN(n688) );
  CLKBUF_X1 U914 ( .A(n1266), .Z(n689) );
  NAND4_X1 U915 ( .A1(n1269), .A2(n1266), .A3(n687), .A4(n633), .ZN(n1253) );
  NOR2_X1 U916 ( .A1(n472), .A2(n1205), .ZN(n691) );
  OR4_X2 U917 ( .A1(n962), .A2(n227), .A3(n965), .A4(n967), .ZN(n974) );
  INV_X1 U918 ( .A(n1299), .ZN(n692) );
  CLKBUF_X1 U919 ( .A(n637), .Z(n693) );
  CLKBUF_X1 U920 ( .A(n1220), .Z(n694) );
  INV_X1 U921 ( .A(n365), .ZN(n695) );
  INV_X1 U922 ( .A(n726), .ZN(n1152) );
  NOR2_X1 U923 ( .A1(n1517), .A2(n82), .ZN(n766) );
  NOR2_X1 U924 ( .A1(n1521), .A2(n728), .ZN(n726) );
  OAI22_X1 U925 ( .A1(n520), .A2(n1678), .B1(n23), .B2(n1896), .ZN(n1892) );
  NAND2_X1 U926 ( .A1(n738), .A2(n696), .ZN(n995) );
  AND2_X1 U927 ( .A1(n988), .A2(n985), .ZN(n696) );
  AND2_X1 U928 ( .A1(n738), .A2(n988), .ZN(n697) );
  NOR2_X1 U929 ( .A1(n689), .A2(n248), .ZN(n699) );
  AND2_X1 U930 ( .A1(n272), .A2(n689), .ZN(n700) );
  NAND2_X1 U931 ( .A1(n1135), .A2(n624), .ZN(n701) );
  NOR2_X1 U932 ( .A1(n702), .A2(n1159), .ZN(n1188) );
  OR2_X1 U933 ( .A1(n1164), .A2(n1163), .ZN(n702) );
  OR2_X1 U934 ( .A1(n873), .A2(n527), .ZN(n869) );
  OR2_X1 U935 ( .A1(n868), .A2(n867), .ZN(n706) );
  NOR2_X1 U936 ( .A1(n1393), .A2(n711), .ZN(n708) );
  NAND2_X1 U937 ( .A1(n391), .A2(n1226), .ZN(n711) );
  OR2_X1 U938 ( .A1(n529), .A2(n1089), .ZN(n1119) );
  AND2_X1 U939 ( .A1(n189), .A2(n239), .ZN(n712) );
  NOR2_X1 U940 ( .A1(n927), .A2(n144), .ZN(n714) );
  NAND2_X1 U941 ( .A1(n734), .A2(n892), .ZN(n715) );
  OR2_X1 U942 ( .A1(n680), .A2(n1074), .ZN(n716) );
  NAND2_X1 U943 ( .A1(n865), .A2(n486), .ZN(n719) );
  NAND2_X1 U944 ( .A1(n718), .A2(n864), .ZN(n720) );
  INV_X1 U945 ( .A(n865), .ZN(n718) );
  XNOR2_X1 U946 ( .A(n960), .B(n649), .ZN(n991) );
  XNOR2_X1 U947 ( .A(n721), .B(n1374), .ZN(n1407) );
  NOR2_X1 U948 ( .A1(n376), .A2(n731), .ZN(n721) );
  NAND2_X1 U949 ( .A1(n1095), .A2(n154), .ZN(n722) );
  NOR2_X1 U950 ( .A1(n1173), .A2(n1174), .ZN(n723) );
  OR2_X1 U951 ( .A1(n1121), .A2(n1118), .ZN(n728) );
  INV_X1 U952 ( .A(n1087), .ZN(n729) );
  NAND2_X1 U953 ( .A1(n567), .A2(n1365), .ZN(n731) );
  NOR2_X1 U954 ( .A1(n1121), .A2(n648), .ZN(n732) );
  AND2_X1 U955 ( .A1(n542), .A2(n781), .ZN(n733) );
  INV_X1 U956 ( .A(n437), .ZN(n894) );
  AOI21_X1 U957 ( .B1(n284), .B2(n626), .A(n736), .ZN(n735) );
  NOR2_X1 U958 ( .A1(n284), .A2(n763), .ZN(n736) );
  OR2_X1 U959 ( .A1(n648), .A2(n1121), .ZN(n1170) );
  OR2_X1 U960 ( .A1(n1903), .A2(n481), .ZN(n1906) );
  AND2_X1 U961 ( .A1(n617), .A2(n1415), .ZN(n737) );
  AND2_X1 U962 ( .A1(n225), .A2(n837), .ZN(n739) );
  AND2_X1 U963 ( .A1(n345), .A2(n179), .ZN(n741) );
  OR2_X1 U964 ( .A1(n1286), .A2(n1287), .ZN(n745) );
  OR2_X1 U965 ( .A1(n120), .A2(n235), .ZN(n1319) );
  INV_X1 U966 ( .A(n434), .ZN(n746) );
  NAND2_X1 U967 ( .A1(n919), .A2(n746), .ZN(n747) );
  CLKBUF_X1 U968 ( .A(n1898), .Z(n748) );
  INV_X1 U969 ( .A(n805), .ZN(n750) );
  INV_X1 U970 ( .A(n750), .ZN(n751) );
  INV_X1 U971 ( .A(n1050), .ZN(n752) );
  INV_X1 U972 ( .A(n630), .ZN(n1050) );
  AOI21_X1 U973 ( .B1(n753), .B2(n1028), .A(n759), .ZN(n758) );
  OR2_X1 U974 ( .A1(n1039), .A2(n284), .ZN(n753) );
  OAI22_X1 U975 ( .A1(n529), .A2(n1555), .B1(n1572), .B2(n147), .ZN(n1782) );
  INV_X1 U976 ( .A(n241), .ZN(n757) );
  NOR2_X1 U977 ( .A1(n763), .A2(n553), .ZN(n759) );
  NOR2_X1 U978 ( .A1(n191), .A2(n251), .ZN(n760) );
  NAND2_X1 U979 ( .A1(n1537), .A2(n1040), .ZN(n763) );
  INV_X1 U980 ( .A(n766), .ZN(n932) );
  INV_X1 U981 ( .A(n883), .ZN(n767) );
  NAND2_X1 U982 ( .A1(n633), .A2(n689), .ZN(n769) );
  NOR2_X1 U983 ( .A1(n425), .A2(n200), .ZN(n771) );
  AND2_X1 U984 ( .A1(n248), .A2(n689), .ZN(n772) );
  NOR2_X1 U985 ( .A1(n773), .A2(n774), .ZN(n782) );
  NOR2_X1 U986 ( .A1(n916), .A2(n652), .ZN(n775) );
  NOR2_X1 U987 ( .A1(n628), .A2(n707), .ZN(n780) );
  NOR2_X1 U988 ( .A1(n49), .A2(n148), .ZN(n785) );
  NOR2_X1 U989 ( .A1(n1668), .A2(n745), .ZN(n776) );
  NAND2_X1 U990 ( .A1(n542), .A2(n117), .ZN(n1071) );
  NOR2_X1 U991 ( .A1(n1050), .A2(n536), .ZN(n781) );
  INV_X1 U992 ( .A(n413), .ZN(n783) );
  NAND3_X1 U993 ( .A1(n588), .A2(n1288), .A3(n1290), .ZN(n1284) );
  NAND3_X1 U994 ( .A1(n688), .A2(n1262), .A3(n1261), .ZN(n1254) );
  AND2_X1 U995 ( .A1(n1367), .A2(n567), .ZN(n786) );
  AND2_X1 U996 ( .A1(n522), .A2(n1190), .ZN(n788) );
  AND2_X1 U997 ( .A1(n185), .A2(n1008), .ZN(n789) );
  OR2_X1 U998 ( .A1(n646), .A2(n1060), .ZN(n1087) );
  OR2_X1 U999 ( .A1(n193), .A2(n200), .ZN(n928) );
  INV_X1 U1000 ( .A(n713), .ZN(n790) );
  NAND3_X1 U1001 ( .A1(n1916), .A2(n1915), .A3(n482), .ZN(n1634) );
  AND2_X2 U1002 ( .A1(n1898), .A2(n96), .ZN(n791) );
  NAND2_X1 U1003 ( .A1(n1401), .A2(n1404), .ZN(n1378) );
  CLKBUF_X1 U1004 ( .A(n1870), .Z(n817) );
  OR2_X1 U1005 ( .A1(n1591), .A2(n824), .ZN(n1549) );
  NAND2_X1 U1006 ( .A1(n1190), .A2(n1192), .ZN(n1173) );
  INV_X1 U1007 ( .A(n643), .ZN(n1589) );
  AOI211_X1 U1008 ( .C1(n96), .C2(n1891), .A(n478), .B(n1890), .ZN(n1632) );
  OR2_X1 U1009 ( .A1(n1581), .A2(n823), .ZN(n1552) );
  INV_X1 U1010 ( .A(n645), .ZN(n1579) );
  CLKBUF_X1 U1011 ( .A(n822), .Z(n812) );
  INV_X1 U1012 ( .A(n151), .ZN(n1569) );
  AOI211_X1 U1013 ( .C1(n438), .C2(n1052), .A(n193), .B(n968), .ZN(n947) );
  INV_X1 U1014 ( .A(a[0]), .ZN(n1918) );
  INV_X1 U1015 ( .A(a[1]), .ZN(n1919) );
  XNOR2_X1 U1016 ( .A(n793), .B(e[3]), .ZN(n834) );
  XNOR2_X1 U1017 ( .A(n794), .B(e[5]), .ZN(n839) );
  XNOR2_X1 U1018 ( .A(n795), .B(e[7]), .ZN(n845) );
  INV_X1 U1019 ( .A(n821), .ZN(n796) );
  BUF_X4 U1020 ( .A(n1526), .Z(n821) );
  AOI211_X1 U1021 ( .C1(n1007), .C2(n1006), .A(n800), .B(n1029), .ZN(n797) );
  AOI211_X1 U1022 ( .C1(n1188), .C2(n1187), .A(n803), .B(n1209), .ZN(n798) );
  OAI21_X1 U1023 ( .B1(n975), .B2(n141), .A(n577), .ZN(n799) );
  OAI21_X1 U1024 ( .B1(n975), .B2(n974), .A(n577), .ZN(n800) );
  CLKBUF_X1 U1025 ( .A(n822), .Z(n811) );
  CLKBUF_X1 U1026 ( .A(n801), .Z(n802) );
  INV_X1 U1027 ( .A(n477), .ZN(n1640) );
  INV_X1 U1028 ( .A(n823), .ZN(n803) );
  INV_X1 U1029 ( .A(n324), .ZN(n1537) );
  AOI211_X1 U1030 ( .C1(n383), .C2(n854), .A(a[22]), .B(n796), .ZN(n807) );
  AOI211_X1 U1031 ( .C1(n111), .C2(n109), .A(n810), .B(n1420), .ZN(n808) );
  NAND4_X1 U1032 ( .A1(n1234), .A2(n1236), .A3(n1238), .A4(n1240), .ZN(n1222)
         );
  OAI21_X1 U1033 ( .B1(n1149), .B2(n1148), .A(n1220), .ZN(n1521) );
  INV_X1 U1034 ( .A(n681), .ZN(n1543) );
  INV_X1 U1035 ( .A(n824), .ZN(n810) );
  OAI21_X1 U1036 ( .B1(n975), .B2(n141), .A(n577), .ZN(n1518) );
  OAI21_X1 U1037 ( .B1(n1437), .B2(n432), .A(n1512), .ZN(n1592) );
  OAI21_X1 U1038 ( .B1(n1038), .B2(n1037), .A(n1081), .ZN(n1183) );
  NAND4_X1 U1039 ( .A1(n79), .A2(n933), .A3(n926), .A4(n929), .ZN(n925) );
  NOR2_X1 U1040 ( .A1(n1378), .A2(n1379), .ZN(n1397) );
  NOR2_X1 U1041 ( .A1(n548), .A2(n72), .ZN(n1398) );
  NOR2_X1 U1042 ( .A1(n1174), .A2(n1173), .ZN(n1187) );
  INV_X1 U1043 ( .A(n1189), .ZN(n1810) );
  NAND4_X1 U1044 ( .A1(n654), .A2(n393), .A3(n1494), .A4(n57), .ZN(n1475) );
  NAND4_X1 U1045 ( .A1(n758), .A2(n1067), .A3(n1072), .A4(n124), .ZN(n1057) );
  NAND4_X1 U1046 ( .A1(n1484), .A2(n1483), .A3(n1480), .A4(n1477), .ZN(n1476)
         );
  NAND4_X1 U1047 ( .A1(n1455), .A2(n1452), .A3(n106), .A4(n1449), .ZN(n1437)
         );
  NAND4_X1 U1048 ( .A1(n621), .A2(n1129), .A3(n624), .A4(n1135), .ZN(n1114) );
  NAND4_X1 U1049 ( .A1(n226), .A2(n964), .A3(n961), .A4(n164), .ZN(n948) );
  INV_X1 U1050 ( .A(n1524), .ZN(n820) );
  NAND4_X1 U1051 ( .A1(n1124), .A2(n1123), .A3(n1120), .A4(n1117), .ZN(n1115)
         );
  XNOR2_X1 U1052 ( .A(n1486), .B(n37), .ZN(n1599) );
  NAND4_X1 U1053 ( .A1(n189), .A2(n78), .A3(n1329), .A4(n1335), .ZN(n1314) );
  NAND4_X1 U1054 ( .A1(n1099), .A2(n1095), .A3(n602), .A4(n1102), .ZN(n1083)
         );
  NAND4_X1 U1055 ( .A1(n1317), .A2(n1320), .A3(n1323), .A4(n1324), .ZN(n1315)
         );
  NAND2_X1 U1056 ( .A1(n1407), .A2(n1408), .ZN(n1379) );
  OAI21_X1 U1057 ( .B1(n60), .B2(n1354), .A(n420), .ZN(n1523) );
  NAND4_X1 U1058 ( .A1(n1368), .A2(n244), .A3(n275), .A4(n1362), .ZN(n1353) );
  NAND4_X1 U1059 ( .A1(n1294), .A2(n287), .A3(n1298), .A4(n698), .ZN(n1283) );
  NAND2_X1 U1060 ( .A1(n1195), .A2(n1194), .ZN(n1174) );
  NAND4_X1 U1061 ( .A1(n1166), .A2(n1171), .A3(n1150), .A4(n1165), .ZN(n1149)
         );
  NAND2_X1 U1062 ( .A1(n862), .A2(n861), .ZN(n852) );
  NOR2_X1 U1063 ( .A1(n852), .A2(n851), .ZN(n854) );
  NAND2_X1 U1064 ( .A1(n1015), .A2(n1016), .ZN(n999) );
  NOR2_X1 U1065 ( .A1(n998), .A2(n999), .ZN(n1006) );
  NAND4_X1 U1066 ( .A1(n1356), .A2(n1376), .A3(n1371), .A4(n75), .ZN(n1354) );
  INV_X1 U1067 ( .A(n820), .ZN(n819) );
  NAND4_X1 U1068 ( .A1(n1599), .A2(n1601), .A3(n1594), .A4(n1597), .ZN(n1515)
         );
  INV_X1 U1069 ( .A(n856), .ZN(n1524) );
  INV_X2 U1070 ( .A(n820), .ZN(n818) );
  INV_X2 U1071 ( .A(n1000), .ZN(n1689) );
  INV_X2 U1072 ( .A(n1001), .ZN(n1687) );
  INV_X2 U1073 ( .A(n1175), .ZN(n1788) );
  INV_X2 U1074 ( .A(n1176), .ZN(n1786) );
  INV_X2 U1075 ( .A(n1380), .ZN(n1856) );
  INV_X2 U1076 ( .A(n1381), .ZN(n1854) );
  INV_X2 U1077 ( .A(n1642), .ZN(n1888) );
  INV_X2 U1078 ( .A(n1643), .ZN(n1883) );
  INV_X1 U1079 ( .A(e[0]), .ZN(n826) );
  XOR2_X1 U1080 ( .A(n410), .B(n826), .Z(n849) );
  NAND4_X1 U1081 ( .A1(n834), .A2(n837), .A3(n849), .A4(n831), .ZN(n830) );
  NAND4_X1 U1082 ( .A1(n845), .A2(n844), .A3(n839), .A4(n842), .ZN(n829) );
  INV_X1 U1083 ( .A(a[23]), .ZN(n876) );
  OAI21_X1 U1084 ( .B1(n829), .B2(n830), .A(n876), .ZN(n853) );
  INV_X1 U1085 ( .A(n414), .ZN(n1526) );
  NOR2_X1 U1086 ( .A1(n1918), .A2(n821), .ZN(normResult[0]) );
  NAND2_X1 U1087 ( .A1(n1526), .A2(n849), .ZN(n848) );
  OAI21_X1 U1088 ( .B1(n831), .B2(n524), .A(n833), .ZN(n832) );
  INV_X1 U1089 ( .A(n832), .ZN(n857) );
  NAND2_X1 U1090 ( .A1(n225), .A2(n837), .ZN(n836) );
  INV_X1 U1091 ( .A(n495), .ZN(n871) );
  OAI21_X1 U1092 ( .B1(n837), .B2(n225), .A(n836), .ZN(n838) );
  INV_X1 U1093 ( .A(n838), .ZN(n874) );
  NAND2_X1 U1094 ( .A1(n618), .A2(n362), .ZN(n841) );
  OAI21_X1 U1095 ( .B1(n216), .B2(n740), .A(n374), .ZN(n840) );
  INV_X1 U1096 ( .A(n840), .ZN(n866) );
  OAI21_X1 U1097 ( .B1(n362), .B2(n618), .A(n841), .ZN(n843) );
  INV_X1 U1098 ( .A(n844), .ZN(n846) );
  OAI21_X1 U1099 ( .B1(n374), .B2(n846), .A(n6), .ZN(n862) );
  OAI21_X1 U1100 ( .B1(n849), .B2(n1526), .A(n848), .ZN(n850) );
  INV_X1 U1101 ( .A(n850), .ZN(n859) );
  NAND2_X1 U1102 ( .A1(n807), .A2(n859), .ZN(n858) );
  OAI21_X1 U1103 ( .B1(n856), .B2(n859), .A(n858), .ZN(n860) );
  INV_X1 U1104 ( .A(n860), .ZN(n881) );
  INV_X1 U1105 ( .A(n873), .ZN(n870) );
  NAND2_X1 U1106 ( .A1(n471), .A2(n485), .ZN(n865) );
  INV_X1 U1107 ( .A(n486), .ZN(n864) );
  INV_X1 U1108 ( .A(n862), .ZN(n863) );
  OAI21_X1 U1109 ( .B1(n864), .B2(n865), .A(n863), .ZN(n884) );
  OAI21_X1 U1110 ( .B1(n373), .B2(n866), .A(n865), .ZN(n867) );
  INV_X1 U1111 ( .A(n334), .ZN(n886) );
  INV_X1 U1112 ( .A(n335), .ZN(n889) );
  OAI21_X1 U1113 ( .B1(n871), .B2(n870), .A(n869), .ZN(n872) );
  INV_X1 U1114 ( .A(n872), .ZN(n892) );
  OAI21_X1 U1115 ( .B1(n874), .B2(n508), .A(n873), .ZN(n875) );
  INV_X1 U1116 ( .A(n875), .ZN(n895) );
  INV_X1 U1117 ( .A(a[22]), .ZN(n897) );
  NAND2_X1 U1118 ( .A1(n1524), .A2(n821), .ZN(n1527) );
  INV_X1 U1119 ( .A(a[21]), .ZN(n921) );
  OAI221_X1 U1120 ( .B1(n897), .B2(n1527), .C1(n819), .C2(n921), .A(n876), 
        .ZN(n877) );
  INV_X1 U1121 ( .A(n877), .ZN(n922) );
  NAND2_X1 U1122 ( .A1(n367), .A2(n881), .ZN(n880) );
  INV_X1 U1123 ( .A(n880), .ZN(n878) );
  OAI21_X1 U1124 ( .B1(n878), .B2(n332), .A(n883), .ZN(n879) );
  INV_X1 U1125 ( .A(n879), .ZN(n901) );
  OAI21_X1 U1126 ( .B1(n881), .B2(n398), .A(n880), .ZN(n882) );
  INV_X1 U1127 ( .A(n484), .ZN(n904) );
  INV_X1 U1128 ( .A(n884), .ZN(n885) );
  OAI21_X1 U1129 ( .B1(n675), .B2(n136), .A(n885), .ZN(n908) );
  XOR2_X1 U1130 ( .A(n515), .B(n675), .Z(n907) );
  OAI21_X1 U1131 ( .B1(n516), .B2(n886), .A(n136), .ZN(n887) );
  INV_X1 U1132 ( .A(n887), .ZN(n911) );
  OAI21_X1 U1133 ( .B1(n445), .B2(n889), .A(n888), .ZN(n890) );
  INV_X1 U1134 ( .A(n890), .ZN(n914) );
  OAI21_X1 U1135 ( .B1(n895), .B2(n767), .A(n894), .ZN(n896) );
  INV_X1 U1136 ( .A(n389), .ZN(n919) );
  INV_X1 U1137 ( .A(a[20]), .ZN(n945) );
  OAI222_X1 U1138 ( .A1(n813), .A2(n921), .B1(n821), .B2(n897), .C1(n818), 
        .C2(n945), .ZN(n1003) );
  INV_X1 U1139 ( .A(n1003), .ZN(n946) );
  INV_X1 U1140 ( .A(n381), .ZN(n1528) );
  INV_X1 U1141 ( .A(n903), .ZN(n900) );
  OAI21_X1 U1142 ( .B1(n900), .B2(n901), .A(n906), .ZN(n902) );
  INV_X1 U1143 ( .A(n902), .ZN(n926) );
  OAI21_X1 U1144 ( .B1(n904), .B2(n1528), .A(n903), .ZN(n905) );
  INV_X1 U1145 ( .A(n905), .ZN(n929) );
  INV_X1 U1146 ( .A(n916), .ZN(n913) );
  INV_X1 U1147 ( .A(n908), .ZN(n909) );
  OAI21_X1 U1148 ( .B1(n280), .B2(n613), .A(n909), .ZN(n933) );
  OAI21_X1 U1149 ( .B1(n775), .B2(n163), .A(n910), .ZN(n912) );
  INV_X1 U1150 ( .A(n912), .ZN(n937) );
  OAI21_X1 U1151 ( .B1(n400), .B2(n913), .A(n545), .ZN(n915) );
  INV_X1 U1152 ( .A(n915), .ZN(n940) );
  INV_X1 U1153 ( .A(n218), .ZN(n942) );
  OAI21_X1 U1154 ( .B1(n175), .B2(n919), .A(n440), .ZN(n920) );
  INV_X1 U1155 ( .A(n920), .ZN(n943) );
  NAND2_X1 U1156 ( .A1(n804), .A2(n382), .ZN(n1561) );
  INV_X1 U1157 ( .A(a[19]), .ZN(n969) );
  OAI222_X1 U1158 ( .A1(n813), .A2(n945), .B1(n821), .B2(n921), .C1(n818), 
        .C2(n969), .ZN(n1031) );
  INV_X1 U1159 ( .A(n1031), .ZN(n1005) );
  OAI221_X1 U1160 ( .B1(n946), .B2(n1561), .C1(n1005), .C2(n379), .A(n922), 
        .ZN(n923) );
  INV_X1 U1161 ( .A(n923), .ZN(n971) );
  OAI21_X1 U1162 ( .B1(n771), .B2(n926), .A(n932), .ZN(n927) );
  INV_X1 U1163 ( .A(n927), .ZN(n950) );
  INV_X1 U1164 ( .A(n930), .ZN(n953) );
  INV_X1 U1165 ( .A(n79), .ZN(n935) );
  NAND2_X1 U1166 ( .A1(n580), .A2(n940), .ZN(n939) );
  INV_X1 U1167 ( .A(n184), .ZN(n934) );
  OAI21_X1 U1168 ( .B1(n936), .B2(n935), .A(n934), .ZN(n957) );
  OAI21_X1 U1169 ( .B1(n782), .B2(n937), .A(n936), .ZN(n938) );
  INV_X1 U1170 ( .A(n938), .ZN(n961) );
  OAI21_X1 U1171 ( .B1(n940), .B2(n580), .A(n939), .ZN(n941) );
  INV_X1 U1172 ( .A(n941), .ZN(n964) );
  OAI21_X1 U1173 ( .B1(n943), .B2(n766), .A(n165), .ZN(n944) );
  INV_X1 U1174 ( .A(a[18]), .ZN(n1002) );
  OAI222_X1 U1175 ( .A1(n813), .A2(n969), .B1(n821), .B2(n945), .C1(n818), 
        .C2(n1002), .ZN(n1052) );
  OAI22_X1 U1176 ( .A1(n1561), .A2(n1005), .B1(n804), .B2(n946), .ZN(n968) );
  INV_X1 U1177 ( .A(n665), .ZN(n1564) );
  NAND2_X1 U1178 ( .A1(n228), .A2(n950), .ZN(n955) );
  OAI21_X1 U1179 ( .B1(n394), .B2(n950), .A(n955), .ZN(n951) );
  INV_X1 U1180 ( .A(n951), .ZN(n976) );
  INV_X1 U1181 ( .A(n954), .ZN(n996) );
  INV_X1 U1182 ( .A(n649), .ZN(n959) );
  INV_X1 U1183 ( .A(n957), .ZN(n958) );
  OAI21_X1 U1184 ( .B1(n959), .B2(n960), .A(n958), .ZN(n992) );
  INV_X1 U1185 ( .A(n962), .ZN(n985) );
  OAI21_X1 U1186 ( .B1(n187), .B2(n179), .A(n963), .ZN(n965) );
  INV_X1 U1187 ( .A(n965), .ZN(n988) );
  INV_X1 U1188 ( .A(n188), .ZN(n979) );
  OAI21_X1 U1189 ( .B1(n130), .B2(n611), .A(n213), .ZN(n967) );
  INV_X1 U1190 ( .A(n533), .ZN(n982) );
  INV_X1 U1191 ( .A(n968), .ZN(n972) );
  NAND2_X1 U1192 ( .A1(n665), .A2(n158), .ZN(n1562) );
  INV_X1 U1193 ( .A(a[17]), .ZN(n1030) );
  OAI222_X1 U1194 ( .A1(n813), .A2(n1002), .B1(n821), .B2(n969), .C1(n818), 
        .C2(n1030), .ZN(n1076) );
  AOI22_X1 U1195 ( .A1(n197), .A2(n1076), .B1(n1683), .B2(n1052), .ZN(n970) );
  OAI211_X1 U1196 ( .C1(n972), .C2(n199), .A(n970), .B(n971), .ZN(n973) );
  INV_X1 U1197 ( .A(n973), .ZN(n1035) );
  INV_X1 U1198 ( .A(n799), .ZN(n1720) );
  INV_X1 U1199 ( .A(n977), .ZN(n1009) );
  INV_X1 U1200 ( .A(n981), .ZN(n978) );
  INV_X1 U1201 ( .A(n535), .ZN(n1024) );
  OAI21_X1 U1202 ( .B1(n982), .B2(n496), .A(n981), .ZN(n983) );
  INV_X1 U1203 ( .A(n531), .ZN(n1027) );
  NAND2_X1 U1204 ( .A1(n390), .A2(n988), .ZN(n987) );
  OAI21_X1 U1205 ( .B1(n697), .B2(n985), .A(n995), .ZN(n986) );
  INV_X1 U1206 ( .A(n562), .ZN(n1019) );
  OAI21_X1 U1207 ( .B1(n390), .B2(n988), .A(n987), .ZN(n989) );
  INV_X1 U1208 ( .A(n989), .ZN(n1021) );
  INV_X1 U1209 ( .A(n638), .ZN(n994) );
  INV_X1 U1210 ( .A(n992), .ZN(n993) );
  OAI21_X1 U1211 ( .B1(n994), .B2(n167), .A(n993), .ZN(n1016) );
  OAI21_X1 U1212 ( .B1(n996), .B2(n1720), .A(n653), .ZN(n997) );
  INV_X1 U1213 ( .A(n192), .ZN(n1012) );
  OAI22_X1 U1214 ( .A1(n804), .A2(n1562), .B1(n85), .B2(n158), .ZN(n1000) );
  INV_X1 U1215 ( .A(n1052), .ZN(n1033) );
  NAND2_X1 U1216 ( .A1(n438), .A2(n98), .ZN(n1644) );
  OAI21_X1 U1217 ( .B1(n85), .B2(n199), .A(n1644), .ZN(n1001) );
  INV_X1 U1218 ( .A(a[16]), .ZN(n1051) );
  OAI222_X1 U1219 ( .A1(n813), .A2(n1030), .B1(n821), .B2(n1002), .C1(n818), 
        .C2(n1051), .ZN(n1107) );
  NAND2_X1 U1220 ( .A1(n98), .A2(n399), .ZN(n1567) );
  OAI221_X1 U1221 ( .B1(n1005), .B2(n1689), .C1(n1033), .C2(n1687), .A(n1004), 
        .ZN(n1029) );
  NAND2_X1 U1222 ( .A1(n797), .A2(n1012), .ZN(n1011) );
  OAI21_X1 U1223 ( .B1(n1012), .B2(n797), .A(n1011), .ZN(n1013) );
  INV_X1 U1224 ( .A(n1013), .ZN(n1040) );
  INV_X1 U1225 ( .A(n1026), .ZN(n1023) );
  INV_X1 U1226 ( .A(n453), .ZN(n1018) );
  INV_X1 U1227 ( .A(n1016), .ZN(n1017) );
  OAI21_X1 U1228 ( .B1(n1018), .B2(n279), .A(n1017), .ZN(n1043) );
  OAI21_X1 U1229 ( .B1(n1021), .B2(n557), .A(n1020), .ZN(n1022) );
  OAI21_X1 U1230 ( .B1(n1023), .B2(n1024), .A(n127), .ZN(n1025) );
  INV_X1 U1231 ( .A(n1029), .ZN(n1056) );
  NAND2_X1 U1232 ( .A1(n822), .A2(n1721), .ZN(n1723) );
  INV_X1 U1233 ( .A(n1076), .ZN(n1054) );
  INV_X1 U1234 ( .A(a[15]), .ZN(n1075) );
  OAI222_X1 U1235 ( .A1(n813), .A2(n1051), .B1(n821), .B2(n1030), .C1(n818), 
        .C2(n1075), .ZN(n1139) );
  AOI222_X1 U1236 ( .A1(n1107), .A2(n695), .B1(n198), .B2(n1139), .C1(n1681), 
        .C2(n1031), .ZN(n1032) );
  OAI221_X1 U1237 ( .B1(n1033), .B2(n1689), .C1(n1054), .C2(n1687), .A(n1032), 
        .ZN(n1034) );
  INV_X1 U1238 ( .A(n1034), .ZN(n1080) );
  OAI221_X1 U1239 ( .B1(n1056), .B2(n1723), .C1(n1080), .C2(n1721), .A(n577), 
        .ZN(n1036) );
  INV_X1 U1240 ( .A(n1036), .ZN(n1081) );
  NAND2_X1 U1241 ( .A1(n1537), .A2(n1040), .ZN(n1039) );
  OAI21_X1 U1242 ( .B1(n308), .B2(n1040), .A(n1039), .ZN(n1041) );
  INV_X1 U1243 ( .A(n162), .ZN(n1059) );
  INV_X1 U1244 ( .A(n380), .ZN(n1045) );
  INV_X1 U1245 ( .A(n1043), .ZN(n1044) );
  OAI21_X1 U1246 ( .B1(n1046), .B2(n1045), .A(n1044), .ZN(n1063) );
  OAI21_X1 U1247 ( .B1(n760), .B2(n241), .A(n388), .ZN(n1047) );
  INV_X1 U1248 ( .A(n1047), .ZN(n1067) );
  OAI21_X1 U1249 ( .B1(n764), .B2(n19), .A(n1048), .ZN(n1049) );
  INV_X1 U1250 ( .A(n1049), .ZN(n1072) );
  INV_X1 U1251 ( .A(n1107), .ZN(n1078) );
  INV_X1 U1252 ( .A(a[14]), .ZN(n1106) );
  OAI222_X1 U1253 ( .A1(n813), .A2(n1075), .B1(n821), .B2(n1051), .C1(n818), 
        .C2(n1106), .ZN(n1178) );
  AOI222_X1 U1254 ( .A1(n1139), .A2(n695), .B1(n198), .B2(n1178), .C1(n1681), 
        .C2(n1052), .ZN(n1053) );
  OAI221_X1 U1255 ( .B1(n1054), .B2(n1689), .C1(n1078), .C2(n1687), .A(n1053), 
        .ZN(n1055) );
  INV_X1 U1256 ( .A(n1055), .ZN(n1111) );
  OAI222_X1 U1257 ( .A1(n811), .A2(n1056), .B1(n1111), .B2(n246), .C1(n1080), 
        .C2(n814), .ZN(n1184) );
  INV_X1 U1258 ( .A(n1184), .ZN(n1112) );
  INV_X1 U1259 ( .A(n140), .ZN(n1534) );
  NAND2_X1 U1260 ( .A1(n411), .A2(n755), .ZN(n1061) );
  OAI21_X1 U1261 ( .B1(n755), .B2(n713), .A(n1061), .ZN(n1058) );
  INV_X1 U1262 ( .A(n1058), .ZN(n1085) );
  OAI21_X1 U1263 ( .B1(n1534), .B2(n1059), .A(n790), .ZN(n1060) );
  INV_X1 U1264 ( .A(n1060), .ZN(n1088) );
  INV_X1 U1265 ( .A(n1069), .ZN(n1066) );
  XOR2_X1 U1266 ( .A(n342), .B(n659), .Z(n1090) );
  INV_X1 U1267 ( .A(n1063), .ZN(n1064) );
  OAI21_X1 U1268 ( .B1(n659), .B2(n1065), .A(n1064), .ZN(n1092) );
  OAI21_X1 U1269 ( .B1(n142), .B2(n1066), .A(n1065), .ZN(n1068) );
  INV_X1 U1270 ( .A(n1068), .ZN(n1095) );
  INV_X1 U1271 ( .A(n1070), .ZN(n1099) );
  OAI21_X1 U1272 ( .B1(n343), .B2(n155), .A(n1071), .ZN(n1073) );
  INV_X1 U1273 ( .A(n1073), .ZN(n1102) );
  INV_X1 U1274 ( .A(n1139), .ZN(n1109) );
  INV_X1 U1275 ( .A(a[13]), .ZN(n1138) );
  OAI222_X1 U1276 ( .A1(n813), .A2(n1106), .B1(n821), .B2(n1075), .C1(n818), 
        .C2(n1138), .ZN(n1211) );
  AOI222_X1 U1277 ( .A1(n1178), .A2(n695), .B1(n198), .B2(n1211), .C1(n1681), 
        .C2(n1076), .ZN(n1077) );
  OAI221_X1 U1278 ( .B1(n1078), .B2(n1689), .C1(n1687), .C2(n1109), .A(n1077), 
        .ZN(n1079) );
  INV_X1 U1279 ( .A(n1079), .ZN(n1143) );
  OAI222_X1 U1280 ( .A1(n1111), .A2(n814), .B1(n1143), .B2(n246), .C1(n812), 
        .C2(n1080), .ZN(n1216) );
  INV_X1 U1281 ( .A(n1216), .ZN(n1186) );
  OAI221_X1 U1282 ( .B1(n1112), .B2(n1555), .C1(n1186), .C2(n644), .A(n1081), 
        .ZN(n1082) );
  INV_X1 U1283 ( .A(n1082), .ZN(n1145) );
  OAI21_X1 U1284 ( .B1(n729), .B2(n1085), .A(n554), .ZN(n1086) );
  INV_X1 U1285 ( .A(n1086), .ZN(n1117) );
  OAI21_X1 U1286 ( .B1(n1088), .B2(n1579), .A(n1087), .ZN(n1089) );
  INV_X1 U1287 ( .A(n1089), .ZN(n1120) );
  INV_X1 U1288 ( .A(n339), .ZN(n1094) );
  INV_X1 U1289 ( .A(n554), .ZN(n1104) );
  NAND2_X1 U1290 ( .A1(n1104), .A2(n278), .ZN(n1103) );
  INV_X1 U1291 ( .A(n707), .ZN(n1098) );
  INV_X1 U1292 ( .A(n1092), .ZN(n1093) );
  OAI21_X1 U1293 ( .B1(n555), .B2(n1094), .A(n1093), .ZN(n1124) );
  OAI21_X1 U1294 ( .B1(n1095), .B2(n780), .A(n555), .ZN(n1096) );
  OAI21_X1 U1295 ( .B1(n154), .B2(n1098), .A(n1097), .ZN(n1100) );
  INV_X1 U1296 ( .A(n1100), .ZN(n1129) );
  OAI21_X1 U1297 ( .B1(n278), .B2(n1104), .A(n1103), .ZN(n1105) );
  INV_X1 U1298 ( .A(n1105), .ZN(n1135) );
  INV_X1 U1299 ( .A(n1178), .ZN(n1141) );
  INV_X1 U1300 ( .A(a[12]), .ZN(n1177) );
  OAI222_X1 U1301 ( .A1(n813), .A2(n1138), .B1(n821), .B2(n1106), .C1(n818), 
        .C2(n1177), .ZN(n1243) );
  AOI222_X1 U1302 ( .A1(n1211), .A2(n695), .B1(n198), .B2(n1243), .C1(n1681), 
        .C2(n1107), .ZN(n1108) );
  OAI221_X1 U1303 ( .B1(n1689), .B2(n1109), .C1(n1687), .C2(n1141), .A(n1108), 
        .ZN(n1110) );
  INV_X1 U1304 ( .A(n1110), .ZN(n1182) );
  OAI222_X1 U1305 ( .A1(n1143), .A2(n814), .B1(n1182), .B2(n246), .C1(n812), 
        .C2(n1111), .ZN(n1248) );
  OAI22_X1 U1306 ( .A1(n1555), .A2(n1186), .B1(n805), .B2(n1112), .ZN(n1137)
         );
  INV_X1 U1307 ( .A(n1659), .ZN(n1574) );
  INV_X1 U1308 ( .A(n1119), .ZN(n1116) );
  OAI21_X1 U1309 ( .B1(n1117), .B2(n1116), .A(n1122), .ZN(n1118) );
  INV_X1 U1310 ( .A(n1118), .ZN(n1150) );
  OAI21_X1 U1311 ( .B1(n1120), .B2(n1574), .A(n663), .ZN(n1121) );
  INV_X1 U1312 ( .A(n1121), .ZN(n1171) );
  INV_X1 U1313 ( .A(n1122), .ZN(n1134) );
  INV_X1 U1314 ( .A(n629), .ZN(n1126) );
  INV_X1 U1315 ( .A(n1124), .ZN(n1125) );
  OAI21_X1 U1316 ( .B1(n1126), .B2(n669), .A(n1125), .ZN(n1166) );
  INV_X1 U1317 ( .A(n1127), .ZN(n1158) );
  OAI21_X1 U1318 ( .B1(n625), .B2(n363), .A(n1128), .ZN(n1130) );
  INV_X1 U1319 ( .A(n1130), .ZN(n1162) );
  OAI21_X1 U1320 ( .B1(n624), .B2(n661), .A(n1131), .ZN(n1132) );
  INV_X1 U1321 ( .A(n1132), .ZN(n1153) );
  OAI21_X1 U1322 ( .B1(n1135), .B2(n1134), .A(n1133), .ZN(n1136) );
  INV_X1 U1323 ( .A(n1136), .ZN(n1155) );
  INV_X1 U1324 ( .A(n1137), .ZN(n1146) );
  NAND2_X1 U1325 ( .A1(n529), .A2(n1579), .ZN(n1572) );
  INV_X1 U1326 ( .A(n1211), .ZN(n1180) );
  INV_X1 U1327 ( .A(a[11]), .ZN(n1210) );
  OAI222_X1 U1328 ( .A1(n813), .A2(n1177), .B1(n821), .B2(n1138), .C1(n818), 
        .C2(n1210), .ZN(n1272) );
  AOI222_X1 U1329 ( .A1(n1243), .A2(n695), .B1(n198), .B2(n1272), .C1(n1681), 
        .C2(n1139), .ZN(n1140) );
  OAI221_X1 U1330 ( .B1(n1689), .B2(n1141), .C1(n1687), .C2(n1180), .A(n1140), 
        .ZN(n1142) );
  INV_X1 U1331 ( .A(n1142), .ZN(n1215) );
  OAI222_X1 U1332 ( .A1(n1182), .A2(n814), .B1(n1215), .B2(n246), .C1(n812), 
        .C2(n1143), .ZN(n1277) );
  AOI22_X1 U1333 ( .A1(n792), .A2(n1277), .B1(n1782), .B2(n1248), .ZN(n1144)
         );
  OAI211_X1 U1334 ( .C1(n1146), .C2(n1572), .A(n1144), .B(n1145), .ZN(n1147)
         );
  INV_X1 U1335 ( .A(n1147), .ZN(n1220) );
  INV_X1 U1336 ( .A(n648), .ZN(n1809) );
  OAI21_X1 U1337 ( .B1(n1150), .B2(n732), .A(n1152), .ZN(n1151) );
  INV_X1 U1338 ( .A(n1151), .ZN(n1190) );
  OAI21_X1 U1339 ( .B1(n601), .B2(n1153), .A(n1157), .ZN(n1154) );
  INV_X1 U1340 ( .A(n325), .ZN(n1204) );
  INV_X1 U1341 ( .A(n1156), .ZN(n1207) );
  INV_X1 U1342 ( .A(n1157), .ZN(n1161) );
  NAND2_X1 U1343 ( .A1(n510), .A2(n1162), .ZN(n1160) );
  OAI21_X1 U1344 ( .B1(n511), .B2(n1158), .A(n513), .ZN(n1159) );
  INV_X1 U1345 ( .A(n571), .ZN(n1199) );
  OAI21_X1 U1346 ( .B1(n1161), .B2(n1162), .A(n1160), .ZN(n1163) );
  INV_X1 U1347 ( .A(n296), .ZN(n1202) );
  INV_X1 U1348 ( .A(n1165), .ZN(n1168) );
  INV_X1 U1349 ( .A(n1166), .ZN(n1167) );
  OAI21_X1 U1350 ( .B1(n1168), .B2(n513), .A(n1167), .ZN(n1195) );
  OAI21_X1 U1351 ( .B1(n1171), .B2(n1809), .A(n1170), .ZN(n1172) );
  INV_X1 U1352 ( .A(n1172), .ZN(n1192) );
  OAI22_X1 U1353 ( .A1(n751), .A2(n1572), .B1(n1555), .B2(n1579), .ZN(n1175)
         );
  INV_X1 U1354 ( .A(n1248), .ZN(n1218) );
  NAND2_X1 U1355 ( .A1(n1534), .A2(n646), .ZN(n1654) );
  OAI21_X1 U1356 ( .B1(n1555), .B2(n1572), .A(n1654), .ZN(n1176) );
  INV_X1 U1357 ( .A(n1243), .ZN(n1213) );
  INV_X1 U1358 ( .A(a[10]), .ZN(n1242) );
  OAI222_X1 U1359 ( .A1(n813), .A2(n1210), .B1(n821), .B2(n1177), .C1(n818), 
        .C2(n1242), .ZN(n1302) );
  AOI222_X1 U1360 ( .A1(n1272), .A2(n695), .B1(n198), .B2(n1302), .C1(n1681), 
        .C2(n1178), .ZN(n1179) );
  OAI221_X1 U1361 ( .B1(n1689), .B2(n1180), .C1(n1687), .C2(n1213), .A(n1179), 
        .ZN(n1181) );
  INV_X1 U1362 ( .A(n1181), .ZN(n1247) );
  OAI222_X1 U1363 ( .A1(n1215), .A2(n814), .B1(n1247), .B2(n246), .C1(n812), 
        .C2(n1182), .ZN(n1307) );
  NAND2_X1 U1364 ( .A1(n645), .A2(n750), .ZN(n1577) );
  OAI221_X1 U1365 ( .B1(n1186), .B2(n1788), .C1(n1218), .C2(n1786), .A(n1185), 
        .ZN(n1209) );
  NAND2_X1 U1366 ( .A1(n3), .A2(n1192), .ZN(n1191) );
  OAI21_X1 U1367 ( .B1(n1192), .B2(n1189), .A(n1191), .ZN(n1193) );
  INV_X1 U1368 ( .A(n1193), .ZN(n1226) );
  NAND2_X1 U1369 ( .A1(n672), .A2(n574), .ZN(n1203) );
  INV_X1 U1370 ( .A(n1194), .ZN(n1197) );
  XOR2_X1 U1371 ( .A(n1198), .B(n1197), .Z(n1228) );
  INV_X1 U1372 ( .A(n1195), .ZN(n1196) );
  OAI21_X1 U1373 ( .B1(n1197), .B2(n214), .A(n1196), .ZN(n1230) );
  OAI21_X1 U1374 ( .B1(n676), .B2(n1199), .A(n214), .ZN(n1200) );
  INV_X1 U1375 ( .A(n1200), .ZN(n1234) );
  INV_X1 U1376 ( .A(n472), .ZN(n1236) );
  OAI21_X1 U1377 ( .B1(n574), .B2(n304), .A(n1203), .ZN(n1205) );
  INV_X1 U1378 ( .A(n1205), .ZN(n1238) );
  OAI21_X1 U1379 ( .B1(n1207), .B2(n788), .A(n1206), .ZN(n1208) );
  INV_X1 U1380 ( .A(n1208), .ZN(n1240) );
  INV_X1 U1381 ( .A(n1209), .ZN(n1252) );
  NAND2_X1 U1382 ( .A1(n1810), .A2(n823), .ZN(n1812) );
  INV_X1 U1383 ( .A(n1277), .ZN(n1250) );
  INV_X1 U1384 ( .A(n1272), .ZN(n1245) );
  INV_X1 U1385 ( .A(a[9]), .ZN(n1271) );
  OAI222_X1 U1386 ( .A1(n813), .A2(n1242), .B1(n821), .B2(n1210), .C1(n818), 
        .C2(n1271), .ZN(n1339) );
  AOI222_X1 U1387 ( .A1(n1302), .A2(n695), .B1(n198), .B2(n1339), .C1(n1681), 
        .C2(n1211), .ZN(n1212) );
  OAI221_X1 U1388 ( .B1(n1689), .B2(n1213), .C1(n1687), .C2(n1245), .A(n1212), 
        .ZN(n1214) );
  INV_X1 U1389 ( .A(n1214), .ZN(n1276) );
  OAI222_X1 U1390 ( .A1(n1247), .A2(n814), .B1(n1276), .B2(n246), .C1(n812), 
        .C2(n1215), .ZN(n1344) );
  AOI222_X1 U1391 ( .A1(n1307), .A2(n679), .B1(n641), .B2(n1344), .C1(n1780), 
        .C2(n1216), .ZN(n1217) );
  OAI221_X1 U1392 ( .B1(n1218), .B2(n1788), .C1(n1250), .C2(n1786), .A(n1217), 
        .ZN(n1219) );
  INV_X1 U1393 ( .A(n1219), .ZN(n1281) );
  OAI221_X1 U1394 ( .B1(n1252), .B2(n1812), .C1(n1281), .C2(n1810), .A(n694), 
        .ZN(n1221) );
  NAND2_X1 U1395 ( .A1(n584), .A2(n572), .ZN(n1229) );
  OAI21_X1 U1396 ( .B1(n572), .B2(n584), .A(n1229), .ZN(n1224) );
  INV_X1 U1397 ( .A(n1224), .ZN(n1255) );
  INV_X1 U1398 ( .A(n1227), .ZN(n1258) );
  INV_X1 U1399 ( .A(n1228), .ZN(n1232) );
  NAND2_X1 U1400 ( .A1(n708), .A2(n1240), .ZN(n1239) );
  INV_X1 U1401 ( .A(n1230), .ZN(n1231) );
  OAI21_X1 U1402 ( .B1(n1232), .B2(n634), .A(n1231), .ZN(n1262) );
  OAI21_X1 U1403 ( .B1(n684), .B2(n581), .A(n1235), .ZN(n1237) );
  INV_X1 U1404 ( .A(n1237), .ZN(n1266) );
  OAI21_X1 U1405 ( .B1(n708), .B2(n1240), .A(n1239), .ZN(n1241) );
  INV_X1 U1406 ( .A(n1241), .ZN(n1269) );
  INV_X1 U1407 ( .A(n1307), .ZN(n1279) );
  INV_X1 U1408 ( .A(n1302), .ZN(n1274) );
  INV_X1 U1409 ( .A(a[8]), .ZN(n1301) );
  OAI222_X1 U1410 ( .A1(n813), .A2(n1271), .B1(n821), .B2(n1242), .C1(n818), 
        .C2(n1301), .ZN(n1383) );
  AOI222_X1 U1411 ( .A1(n1339), .A2(n695), .B1(n198), .B2(n1383), .C1(n1681), 
        .C2(n1243), .ZN(n1244) );
  OAI221_X1 U1412 ( .B1(n1689), .B2(n1245), .C1(n1687), .C2(n1274), .A(n1244), 
        .ZN(n1246) );
  INV_X1 U1413 ( .A(n1246), .ZN(n1306) );
  OAI222_X1 U1414 ( .A1(n1276), .A2(n814), .B1(n1306), .B2(n246), .C1(n812), 
        .C2(n1247), .ZN(n1388) );
  AOI222_X1 U1415 ( .A1(n1344), .A2(n679), .B1(n641), .B2(n1388), .C1(n1780), 
        .C2(n1248), .ZN(n1249) );
  OAI221_X1 U1416 ( .B1(n1250), .B2(n1788), .C1(n1279), .C2(n1786), .A(n1249), 
        .ZN(n1251) );
  INV_X1 U1417 ( .A(n1251), .ZN(n1311) );
  OAI222_X1 U1418 ( .A1(n823), .A2(n1252), .B1(n1311), .B2(n397), .C1(n1281), 
        .C2(n815), .ZN(n1394) );
  INV_X1 U1419 ( .A(n1394), .ZN(n1312) );
  INV_X1 U1420 ( .A(n415), .ZN(n1540) );
  OAI21_X1 U1421 ( .B1(n319), .B2(n1255), .A(n1260), .ZN(n1256) );
  INV_X1 U1422 ( .A(n170), .ZN(n1285) );
  NAND2_X1 U1423 ( .A1(n677), .A2(n402), .ZN(n1268) );
  XOR2_X1 U1424 ( .A(n89), .B(n635), .Z(n1288) );
  INV_X1 U1425 ( .A(n1262), .ZN(n1263) );
  OAI21_X1 U1426 ( .B1(n635), .B2(n1264), .A(n1263), .ZN(n1290) );
  OAI21_X1 U1427 ( .B1(n772), .B2(n633), .A(n89), .ZN(n1265) );
  INV_X1 U1428 ( .A(n1265), .ZN(n1294) );
  OAI21_X1 U1429 ( .B1(n779), .B2(n686), .A(n267), .ZN(n1267) );
  INV_X1 U1430 ( .A(n1267), .ZN(n1298) );
  OAI21_X1 U1431 ( .B1(n402), .B2(n677), .A(n1268), .ZN(n1270) );
  NAND2_X1 U1432 ( .A1(n809), .A2(n415), .ZN(n1551) );
  INV_X1 U1433 ( .A(n1344), .ZN(n1309) );
  INV_X1 U1434 ( .A(n1339), .ZN(n1304) );
  INV_X1 U1435 ( .A(a[7]), .ZN(n1338) );
  OAI222_X1 U1436 ( .A1(n813), .A2(n1301), .B1(n821), .B2(n1271), .C1(n818), 
        .C2(n1338), .ZN(n1422) );
  AOI222_X1 U1437 ( .A1(n1383), .A2(n695), .B1(n198), .B2(n1422), .C1(n1681), 
        .C2(n1272), .ZN(n1273) );
  OAI221_X1 U1438 ( .B1(n1689), .B2(n1274), .C1(n1687), .C2(n1304), .A(n1273), 
        .ZN(n1275) );
  INV_X1 U1439 ( .A(n1275), .ZN(n1343) );
  OAI222_X1 U1440 ( .A1(n1306), .A2(n814), .B1(n1343), .B2(n246), .C1(n812), 
        .C2(n1276), .ZN(n1427) );
  AOI222_X1 U1441 ( .A1(n1388), .A2(n679), .B1(n641), .B2(n1427), .C1(n1780), 
        .C2(n1277), .ZN(n1278) );
  OAI221_X1 U1442 ( .B1(n1279), .B2(n1788), .C1(n1786), .C2(n1309), .A(n1278), 
        .ZN(n1280) );
  INV_X1 U1443 ( .A(n1280), .ZN(n1348) );
  OAI222_X1 U1444 ( .A1(n1311), .A2(n815), .B1(n1348), .B2(n397), .C1(n823), 
        .C2(n1281), .ZN(n1432) );
  INV_X1 U1445 ( .A(n1432), .ZN(n1396) );
  OAI221_X1 U1446 ( .B1(n1312), .B2(n1551), .C1(n1396), .C2(n268), .A(n512), 
        .ZN(n1282) );
  INV_X1 U1447 ( .A(n1282), .ZN(n1350) );
  NAND2_X1 U1448 ( .A1(n639), .A2(n1285), .ZN(n1289) );
  OAI21_X1 U1449 ( .B1(n1285), .B2(n639), .A(n1289), .ZN(n1286) );
  INV_X1 U1450 ( .A(n1286), .ZN(n1317) );
  OAI21_X1 U1451 ( .B1(n221), .B2(n1589), .A(n114), .ZN(n1287) );
  INV_X1 U1452 ( .A(n1287), .ZN(n1320) );
  INV_X1 U1453 ( .A(n210), .ZN(n1292) );
  INV_X1 U1454 ( .A(n1290), .ZN(n1291) );
  OAI21_X1 U1455 ( .B1(n264), .B2(n1292), .A(n1291), .ZN(n1324) );
  OAI21_X1 U1456 ( .B1(n610), .B2(n787), .A(n1293), .ZN(n1295) );
  INV_X1 U1457 ( .A(n1295), .ZN(n1326) );
  OAI21_X1 U1458 ( .B1(n596), .B2(n83), .A(n1296), .ZN(n1297) );
  INV_X1 U1459 ( .A(n1297), .ZN(n1329) );
  OAI21_X1 U1460 ( .B1(n525), .B2(n321), .A(n1299), .ZN(n1300) );
  INV_X1 U1461 ( .A(n1300), .ZN(n1335) );
  INV_X1 U1462 ( .A(n1388), .ZN(n1346) );
  INV_X1 U1463 ( .A(n1383), .ZN(n1341) );
  INV_X1 U1464 ( .A(a[6]), .ZN(n1382) );
  OAI222_X1 U1465 ( .A1(n813), .A2(n1338), .B1(n821), .B2(n1301), .C1(n818), 
        .C2(n1382), .ZN(n1460) );
  AOI222_X1 U1466 ( .A1(n1422), .A2(n695), .B1(n198), .B2(n1460), .C1(n1681), 
        .C2(n1302), .ZN(n1303) );
  OAI221_X1 U1467 ( .B1(n1689), .B2(n1304), .C1(n1687), .C2(n1341), .A(n1303), 
        .ZN(n1305) );
  INV_X1 U1468 ( .A(n1305), .ZN(n1387) );
  OAI222_X1 U1469 ( .A1(n1343), .A2(n814), .B1(n1387), .B2(n246), .C1(n812), 
        .C2(n1306), .ZN(n1465) );
  AOI222_X1 U1470 ( .A1(n1427), .A2(n679), .B1(n641), .B2(n1465), .C1(n1780), 
        .C2(n1307), .ZN(n1308) );
  OAI221_X1 U1471 ( .B1(n1788), .B2(n1309), .C1(n1786), .C2(n1346), .A(n1308), 
        .ZN(n1310) );
  INV_X1 U1472 ( .A(n1310), .ZN(n1392) );
  OAI222_X1 U1473 ( .A1(n1348), .A2(n815), .B1(n1392), .B2(n397), .C1(n823), 
        .C2(n1311), .ZN(n1470) );
  OAI22_X1 U1474 ( .A1(n1551), .A2(n1396), .B1(n809), .B2(n1312), .ZN(n1337)
         );
  INV_X1 U1475 ( .A(n139), .ZN(n1584) );
  INV_X1 U1476 ( .A(n1319), .ZN(n1316) );
  OAI21_X1 U1477 ( .B1(n62), .B2(n1316), .A(n1322), .ZN(n1318) );
  INV_X1 U1478 ( .A(n53), .ZN(n1356) );
  OAI21_X1 U1479 ( .B1(n1584), .B2(n1320), .A(n1319), .ZN(n1321) );
  INV_X1 U1480 ( .A(n1321), .ZN(n1376) );
  INV_X1 U1481 ( .A(n1334), .ZN(n1332) );
  NAND2_X1 U1482 ( .A1(n776), .A2(n712), .ZN(n1331) );
  INV_X1 U1483 ( .A(n1324), .ZN(n1325) );
  OAI21_X1 U1484 ( .B1(n234), .B2(n292), .A(n1325), .ZN(n1372) );
  OAI21_X1 U1485 ( .B1(n293), .B2(n146), .A(n118), .ZN(n1327) );
  INV_X1 U1486 ( .A(n1327), .ZN(n1365) );
  OAI21_X1 U1487 ( .B1(n744), .B2(n323), .A(n1328), .ZN(n1330) );
  INV_X1 U1488 ( .A(n1330), .ZN(n1368) );
  OAI21_X1 U1489 ( .B1(n1332), .B2(n543), .A(n347), .ZN(n1333) );
  INV_X1 U1490 ( .A(n138), .ZN(n1359) );
  OAI21_X1 U1491 ( .B1(n131), .B2(n283), .A(n1334), .ZN(n1336) );
  INV_X1 U1492 ( .A(n1336), .ZN(n1362) );
  INV_X1 U1493 ( .A(n1337), .ZN(n1351) );
  NAND2_X1 U1494 ( .A1(n651), .A2(n1589), .ZN(n1582) );
  INV_X1 U1495 ( .A(n1427), .ZN(n1390) );
  INV_X1 U1496 ( .A(n1422), .ZN(n1385) );
  INV_X1 U1497 ( .A(a[5]), .ZN(n1421) );
  OAI222_X1 U1498 ( .A1(n813), .A2(n1382), .B1(n821), .B2(n1338), .C1(n818), 
        .C2(n1421), .ZN(n1497) );
  AOI222_X1 U1499 ( .A1(n1460), .A2(n695), .B1(n198), .B2(n1497), .C1(n1681), 
        .C2(n1339), .ZN(n1340) );
  OAI221_X1 U1500 ( .B1(n1689), .B2(n1341), .C1(n1687), .C2(n1385), .A(n1340), 
        .ZN(n1342) );
  INV_X1 U1501 ( .A(n1342), .ZN(n1426) );
  OAI222_X1 U1502 ( .A1(n1387), .A2(n814), .B1(n1426), .B2(n246), .C1(n812), 
        .C2(n1343), .ZN(n1502) );
  AOI222_X1 U1503 ( .A1(n1465), .A2(n679), .B1(n641), .B2(n1502), .C1(n1780), 
        .C2(n1344), .ZN(n1345) );
  OAI221_X1 U1504 ( .B1(n1788), .B2(n1346), .C1(n1786), .C2(n1390), .A(n1345), 
        .ZN(n1347) );
  INV_X1 U1505 ( .A(n1347), .ZN(n1431) );
  OAI222_X1 U1506 ( .A1(n1392), .A2(n815), .B1(n1431), .B2(n397), .C1(n823), 
        .C2(n1348), .ZN(n1507) );
  AOI22_X1 U1507 ( .A1(n314), .A2(n1507), .B1(n77), .B2(n1470), .ZN(n1349) );
  OAI211_X1 U1508 ( .C1(n1351), .C2(n350), .A(n1349), .B(n1350), .ZN(n1352) );
  INV_X1 U1509 ( .A(n422), .ZN(n1867) );
  INV_X1 U1510 ( .A(n1375), .ZN(n1355) );
  OAI21_X1 U1511 ( .B1(n1355), .B2(n50), .A(n1358), .ZN(n1357) );
  INV_X1 U1512 ( .A(n1357), .ZN(n1401) );
  NAND2_X1 U1513 ( .A1(n115), .A2(n1359), .ZN(n1364) );
  OAI21_X1 U1514 ( .B1(n657), .B2(n1359), .A(n1364), .ZN(n1360) );
  INV_X1 U1515 ( .A(n316), .ZN(n1418) );
  OAI21_X1 U1516 ( .B1(n1362), .B2(n372), .A(n1361), .ZN(n1363) );
  INV_X1 U1517 ( .A(n87), .ZN(n1419) );
  INV_X1 U1518 ( .A(n1364), .ZN(n1367) );
  INV_X1 U1519 ( .A(n493), .ZN(n1412) );
  OAI21_X1 U1520 ( .B1(n567), .B2(n1367), .A(n1366), .ZN(n1369) );
  INV_X1 U1521 ( .A(n1369), .ZN(n1415) );
  INV_X1 U1522 ( .A(n1371), .ZN(n1374) );
  INV_X1 U1523 ( .A(n76), .ZN(n1373) );
  OAI21_X1 U1524 ( .B1(n724), .B2(n1374), .A(n1373), .ZN(n1408) );
  OAI21_X1 U1525 ( .B1(n1376), .B2(n1867), .A(n1375), .ZN(n1377) );
  INV_X1 U1526 ( .A(n1377), .ZN(n1404) );
  OAI22_X1 U1527 ( .A1(n809), .A2(n1582), .B1(n1551), .B2(n252), .ZN(n1380) );
  INV_X1 U1528 ( .A(n1470), .ZN(n1434) );
  NAND2_X1 U1529 ( .A1(n1540), .A2(n51), .ZN(n1663) );
  OAI21_X1 U1530 ( .B1(n1551), .B2(n350), .A(n1663), .ZN(n1381) );
  INV_X1 U1531 ( .A(n1465), .ZN(n1429) );
  INV_X1 U1532 ( .A(n1460), .ZN(n1424) );
  INV_X1 U1533 ( .A(a[4]), .ZN(n1459) );
  OAI222_X1 U1534 ( .A1(n813), .A2(n1421), .B1(n821), .B2(n1382), .C1(n818), 
        .C2(n1459), .ZN(n1615) );
  AOI222_X1 U1535 ( .A1(n1497), .A2(n695), .B1(n198), .B2(n1615), .C1(n1681), 
        .C2(n1383), .ZN(n1384) );
  OAI221_X1 U1536 ( .B1(n1689), .B2(n1385), .C1(n1687), .C2(n1424), .A(n1384), 
        .ZN(n1386) );
  INV_X1 U1537 ( .A(n1386), .ZN(n1464) );
  OAI222_X1 U1538 ( .A1(n1426), .A2(n814), .B1(n1464), .B2(n246), .C1(n812), 
        .C2(n1387), .ZN(n1621) );
  AOI222_X1 U1539 ( .A1(n1502), .A2(n631), .B1(n641), .B2(n1621), .C1(n1780), 
        .C2(n1388), .ZN(n1389) );
  OAI221_X1 U1540 ( .B1(n1788), .B2(n1390), .C1(n1786), .C2(n1429), .A(n1389), 
        .ZN(n1391) );
  INV_X1 U1541 ( .A(n1391), .ZN(n1469) );
  OAI222_X1 U1542 ( .A1(n1431), .A2(n815), .B1(n1469), .B2(n397), .C1(n823), 
        .C2(n1392), .ZN(n1626) );
  NAND2_X1 U1543 ( .A1(n51), .A2(n682), .ZN(n1587) );
  OAI221_X1 U1544 ( .B1(n1396), .B2(n1856), .C1(n1434), .C2(n1854), .A(n1395), 
        .ZN(n1420) );
  NAND2_X1 U1545 ( .A1(n116), .A2(n1404), .ZN(n1403) );
  INV_X1 U1546 ( .A(n1403), .ZN(n1400) );
  OAI21_X1 U1547 ( .B1(n67), .B2(n1400), .A(n1406), .ZN(n1402) );
  INV_X1 U1548 ( .A(n1402), .ZN(n1438) );
  OAI21_X1 U1549 ( .B1(n1404), .B2(n368), .A(n1403), .ZN(n1405) );
  INV_X1 U1550 ( .A(n1405), .ZN(n1441) );
  NAND2_X1 U1551 ( .A1(n617), .A2(n1415), .ZN(n1414) );
  NAND2_X1 U1552 ( .A1(n637), .A2(n521), .ZN(n1411) );
  INV_X1 U1553 ( .A(n550), .ZN(n1410) );
  INV_X1 U1554 ( .A(n549), .ZN(n1409) );
  OAI21_X1 U1555 ( .B1(n1410), .B2(n1411), .A(n1409), .ZN(n1445) );
  OAI21_X1 U1556 ( .B1(n1412), .B2(n737), .A(n1411), .ZN(n1413) );
  INV_X1 U1557 ( .A(n1413), .ZN(n1449) );
  OAI21_X1 U1558 ( .B1(n1415), .B2(n492), .A(n1414), .ZN(n1416) );
  INV_X1 U1559 ( .A(n1416), .ZN(n1452) );
  INV_X1 U1560 ( .A(n100), .ZN(n1455) );
  INV_X1 U1561 ( .A(n1420), .ZN(n1474) );
  INV_X1 U1562 ( .A(n1507), .ZN(n1472) );
  INV_X1 U1563 ( .A(n1502), .ZN(n1467) );
  INV_X1 U1564 ( .A(n1497), .ZN(n1462) );
  INV_X1 U1565 ( .A(a[3]), .ZN(n1496) );
  OAI222_X1 U1566 ( .A1(n813), .A2(n1459), .B1(n821), .B2(n1421), .C1(n818), 
        .C2(n1496), .ZN(n1680) );
  AOI222_X1 U1567 ( .A1(n1615), .A2(n695), .B1(n198), .B2(n1680), .C1(n1681), 
        .C2(n1422), .ZN(n1423) );
  OAI221_X1 U1568 ( .B1(n1689), .B2(n1424), .C1(n1687), .C2(n1462), .A(n1423), 
        .ZN(n1425) );
  INV_X1 U1569 ( .A(n1425), .ZN(n1501) );
  OAI222_X1 U1570 ( .A1(n1464), .A2(n814), .B1(n1501), .B2(n246), .C1(n812), 
        .C2(n1426), .ZN(n1779) );
  AOI222_X1 U1571 ( .A1(n1621), .A2(n679), .B1(n641), .B2(n1779), .C1(n1780), 
        .C2(n1427), .ZN(n1428) );
  OAI221_X1 U1572 ( .B1(n1788), .B2(n1429), .C1(n1786), .C2(n1467), .A(n1428), 
        .ZN(n1430) );
  INV_X1 U1573 ( .A(n1430), .ZN(n1506) );
  OAI222_X1 U1574 ( .A1(n1469), .A2(n815), .B1(n1506), .B2(n397), .C1(n823), 
        .C2(n1431), .ZN(n1848) );
  AOI222_X1 U1575 ( .A1(n1626), .A2(n730), .B1(n315), .B2(n1848), .C1(n1849), 
        .C2(n1432), .ZN(n1433) );
  OAI221_X1 U1576 ( .B1(n1434), .B2(n1856), .C1(n1472), .C2(n1854), .A(n1433), 
        .ZN(n1435) );
  INV_X1 U1577 ( .A(n1435), .ZN(n1511) );
  OAI221_X1 U1578 ( .B1(n1474), .B2(n816), .C1(n1511), .C2(n1868), .A(n582), 
        .ZN(n1436) );
  INV_X1 U1579 ( .A(n1436), .ZN(n1512) );
  OAI21_X1 U1580 ( .B1(n65), .B2(n636), .A(n1444), .ZN(n1439) );
  INV_X1 U1581 ( .A(n1439), .ZN(n1477) );
  OAI21_X1 U1582 ( .B1(n801), .B2(n1441), .A(n1440), .ZN(n1442) );
  INV_X1 U1583 ( .A(n1442), .ZN(n1480) );
  INV_X1 U1584 ( .A(n1443), .ZN(n1447) );
  INV_X1 U1585 ( .A(n1444), .ZN(n1457) );
  NAND2_X1 U1586 ( .A1(n504), .A2(n500), .ZN(n1454) );
  INV_X1 U1587 ( .A(n149), .ZN(n1451) );
  INV_X1 U1588 ( .A(n1445), .ZN(n1446) );
  OAI21_X1 U1589 ( .B1(n1447), .B2(n674), .A(n1446), .ZN(n1484) );
  OAI21_X1 U1590 ( .B1(n409), .B2(n1449), .A(n674), .ZN(n1450) );
  INV_X1 U1591 ( .A(n309), .ZN(n1487) );
  OAI21_X1 U1592 ( .B1(n1451), .B2(n58), .A(n671), .ZN(n1453) );
  INV_X1 U1593 ( .A(n71), .ZN(n1489) );
  OAI21_X1 U1594 ( .B1(n658), .B2(n488), .A(n149), .ZN(n1456) );
  OAI21_X1 U1595 ( .B1(n1457), .B2(n489), .A(n501), .ZN(n1458) );
  INV_X1 U1596 ( .A(n1458), .ZN(n1494) );
  INV_X1 U1597 ( .A(n1626), .ZN(n1509) );
  INV_X1 U1598 ( .A(n1621), .ZN(n1504) );
  INV_X1 U1599 ( .A(n1615), .ZN(n1499) );
  INV_X1 U1600 ( .A(a[2]), .ZN(n1525) );
  OAI222_X1 U1601 ( .A1(n813), .A2(n1496), .B1(n821), .B2(n1459), .C1(n818), 
        .C2(n1525), .ZN(n1648) );
  AOI222_X1 U1602 ( .A1(n1680), .A2(n695), .B1(n198), .B2(n1648), .C1(n1681), 
        .C2(n1460), .ZN(n1461) );
  OAI221_X1 U1603 ( .B1(n1689), .B2(n1462), .C1(n1687), .C2(n1499), .A(n1461), 
        .ZN(n1463) );
  INV_X1 U1604 ( .A(n1463), .ZN(n1620) );
  OAI222_X1 U1605 ( .A1(n1501), .A2(n814), .B1(n1620), .B2(n246), .C1(n812), 
        .C2(n1464), .ZN(n1765) );
  AOI222_X1 U1606 ( .A1(n1779), .A2(n631), .B1(n641), .B2(n1765), .C1(n1780), 
        .C2(n1465), .ZN(n1466) );
  OAI221_X1 U1607 ( .B1(n1788), .B2(n1467), .C1(n1786), .C2(n1504), .A(n1466), 
        .ZN(n1468) );
  INV_X1 U1608 ( .A(n1468), .ZN(n1625) );
  OAI222_X1 U1609 ( .A1(n1506), .A2(n815), .B1(n1625), .B2(n397), .C1(n823), 
        .C2(n1469), .ZN(n1839) );
  AOI222_X1 U1610 ( .A1(n1848), .A2(n730), .B1(n315), .B2(n1839), .C1(n1849), 
        .C2(n1470), .ZN(n1471) );
  OAI221_X1 U1611 ( .B1(n1472), .B2(n1856), .C1(n1509), .C2(n1854), .A(n1471), 
        .ZN(n1473) );
  INV_X1 U1612 ( .A(n1473), .ZN(n1630) );
  OAI222_X1 U1613 ( .A1(n824), .A2(n1474), .B1(n1630), .B2(n1868), .C1(n1511), 
        .C2(n817), .ZN(n1882) );
  INV_X1 U1614 ( .A(n1882), .ZN(n1631) );
  INV_X1 U1615 ( .A(n312), .ZN(n1679) );
  NAND2_X1 U1616 ( .A1(n36), .A2(n1477), .ZN(n1482) );
  OAI21_X1 U1617 ( .B1(n1477), .B2(n36), .A(n1482), .ZN(n1478) );
  INV_X1 U1618 ( .A(n1478), .ZN(n1594) );
  OAI21_X1 U1619 ( .B1(n1480), .B2(n1679), .A(n1479), .ZN(n1481) );
  INV_X1 U1620 ( .A(n1481), .ZN(n1597) );
  INV_X1 U1621 ( .A(n44), .ZN(n1492) );
  INV_X1 U1622 ( .A(n1484), .ZN(n1485) );
  OAI21_X1 U1623 ( .B1(n1486), .B2(n90), .A(n1485), .ZN(n1601) );
  OAI21_X1 U1624 ( .B1(n1489), .B2(n710), .A(n1488), .ZN(n1490) );
  INV_X1 U1625 ( .A(n39), .ZN(n1608) );
  INV_X1 U1626 ( .A(n41), .ZN(n1611) );
  OAI21_X1 U1627 ( .B1(n785), .B2(n68), .A(n1493), .ZN(n1495) );
  INV_X1 U1628 ( .A(n1495), .ZN(n1614) );
  NAND2_X1 U1629 ( .A1(n46), .A2(n801), .ZN(n1678) );
  INV_X1 U1630 ( .A(n1848), .ZN(n1628) );
  INV_X1 U1631 ( .A(n1779), .ZN(n1623) );
  INV_X1 U1632 ( .A(n1680), .ZN(n1618) );
  OAI222_X1 U1633 ( .A1(n813), .A2(n1525), .B1(n821), .B2(n1496), .C1(n1919), 
        .C2(n818), .ZN(n1616) );
  AOI222_X1 U1634 ( .A1(n1648), .A2(n695), .B1(n198), .B2(n1616), .C1(n1681), 
        .C2(n1497), .ZN(n1498) );
  OAI221_X1 U1635 ( .B1(n1689), .B2(n1499), .C1(n1687), .C2(n1618), .A(n1498), 
        .ZN(n1500) );
  INV_X1 U1636 ( .A(n1500), .ZN(n1719) );
  OAI222_X1 U1637 ( .A1(n1620), .A2(n814), .B1(n1719), .B2(n246), .C1(n812), 
        .C2(n1501), .ZN(n1764) );
  AOI222_X1 U1638 ( .A1(n1765), .A2(n679), .B1(n641), .B2(n1764), .C1(n1780), 
        .C2(n1502), .ZN(n1503) );
  OAI221_X1 U1639 ( .B1(n1788), .B2(n1504), .C1(n1786), .C2(n1623), .A(n1503), 
        .ZN(n1505) );
  INV_X1 U1640 ( .A(n1505), .ZN(n1808) );
  OAI222_X1 U1641 ( .A1(n1625), .A2(n815), .B1(n1808), .B2(n397), .C1(n823), 
        .C2(n1506), .ZN(n1838) );
  AOI222_X1 U1642 ( .A1(n1839), .A2(n730), .B1(n315), .B2(n1838), .C1(n1849), 
        .C2(n1507), .ZN(n1508) );
  OAI221_X1 U1643 ( .B1(n1509), .B2(n1856), .C1(n1854), .C2(n1628), .A(n1508), 
        .ZN(n1510) );
  INV_X1 U1644 ( .A(n1510), .ZN(n1866) );
  OAI222_X1 U1645 ( .A1(n1630), .A2(n817), .B1(n1866), .B2(n366), .C1(n824), 
        .C2(n1511), .ZN(n1878) );
  INV_X1 U1646 ( .A(n1878), .ZN(n1889) );
  OAI221_X1 U1647 ( .B1(n1631), .B2(n1678), .C1(n1889), .C2(n666), .A(n494), 
        .ZN(n1513) );
  INV_X1 U1648 ( .A(n1513), .ZN(n1895) );
  INV_X1 U1649 ( .A(n478), .ZN(n1641) );
  OAI22_X1 U1650 ( .A1(n1918), .A2(n813), .B1(n1919), .B2(n821), .ZN(n1682) );
  NAND2_X1 U1651 ( .A1(n1682), .A2(n399), .ZN(n1529) );
  INV_X1 U1652 ( .A(n1529), .ZN(n1516) );
  NAND2_X1 U1653 ( .A1(n585), .A2(n1516), .ZN(n1532) );
  INV_X1 U1654 ( .A(n1532), .ZN(n1563) );
  NAND2_X1 U1655 ( .A1(n98), .A2(n1563), .ZN(n1571) );
  INV_X1 U1656 ( .A(n1571), .ZN(n1519) );
  NAND2_X1 U1657 ( .A1(n1519), .A2(n799), .ZN(n1556) );
  INV_X1 U1658 ( .A(n1556), .ZN(n1692) );
  NAND2_X1 U1659 ( .A1(n147), .A2(n1692), .ZN(n1538) );
  INV_X1 U1660 ( .A(n1538), .ZN(n1573) );
  NAND2_X1 U1661 ( .A1(n1573), .A2(n645), .ZN(n1581) );
  INV_X1 U1662 ( .A(n1552), .ZN(n1697) );
  NAND2_X1 U1663 ( .A1(n268), .A2(n1697), .ZN(n1544) );
  INV_X1 U1664 ( .A(n1544), .ZN(n1583) );
  NAND2_X1 U1665 ( .A1(n1583), .A2(n51), .ZN(n1591) );
  INV_X1 U1666 ( .A(n1549), .ZN(n1702) );
  NAND2_X1 U1667 ( .A1(n23), .A2(n1702), .ZN(n1635) );
  NOR2_X1 U1668 ( .A1(n1641), .A2(n1635), .ZN(normResult[1]) );
  OAI222_X1 U1669 ( .A1(n1919), .A2(n813), .B1(n821), .B2(n1525), .C1(n1918), 
        .C2(n818), .ZN(n1684) );
  INV_X1 U1670 ( .A(n1684), .ZN(n1560) );
  NAND2_X1 U1671 ( .A1(n804), .A2(n1682), .ZN(n1530) );
  MUX2_X1 U1672 ( .A(n1530), .B(n1529), .S(n438), .Z(n1531) );
  OAI21_X1 U1673 ( .B1(n804), .B2(n1560), .A(n1531), .ZN(n1565) );
  INV_X1 U1674 ( .A(n1565), .ZN(n1651) );
  OAI22_X1 U1675 ( .A1(n1532), .A2(n223), .B1(n158), .B2(n1651), .ZN(n1533) );
  INV_X1 U1676 ( .A(n1533), .ZN(n1653) );
  OAI22_X1 U1677 ( .A1(n814), .A2(n1571), .B1(n812), .B2(n1653), .ZN(n1706) );
  INV_X1 U1678 ( .A(n1706), .ZN(n1554) );
  NAND2_X1 U1679 ( .A1(n1692), .A2(n805), .ZN(n1535) );
  MUX2_X1 U1680 ( .A(n1535), .B(n1556), .S(n1534), .Z(n1536) );
  OAI21_X1 U1681 ( .B1(n751), .B2(n1554), .A(n1536), .ZN(n1575) );
  INV_X1 U1682 ( .A(n1575), .ZN(n1660) );
  OAI22_X1 U1683 ( .A1(n1538), .A2(n619), .B1(n1579), .B2(n1660), .ZN(n1539)
         );
  INV_X1 U1684 ( .A(n1539), .ZN(n1662) );
  OAI22_X1 U1685 ( .A1(n815), .A2(n1581), .B1(n823), .B2(n1662), .ZN(n1711) );
  INV_X1 U1686 ( .A(n1711), .ZN(n1550) );
  NAND2_X1 U1687 ( .A1(n1697), .A2(n809), .ZN(n1541) );
  MUX2_X1 U1688 ( .A(n1541), .B(n1552), .S(n1540), .Z(n1542) );
  OAI21_X1 U1689 ( .B1(n809), .B2(n1550), .A(n1542), .ZN(n1585) );
  INV_X1 U1690 ( .A(n1585), .ZN(n1669) );
  OAI22_X1 U1691 ( .A1(n1544), .A2(n475), .B1(n252), .B2(n1669), .ZN(n1545) );
  INV_X1 U1692 ( .A(n1545), .ZN(n1671) );
  OAI22_X1 U1693 ( .A1(n816), .A2(n1591), .B1(n824), .B2(n1671), .ZN(n1716) );
  INV_X1 U1694 ( .A(n1716), .ZN(n1548) );
  NAND2_X1 U1695 ( .A1(n1702), .A2(n801), .ZN(n1546) );
  MUX2_X1 U1696 ( .A(n1546), .B(n1549), .S(n96), .Z(n1547) );
  OAI21_X1 U1697 ( .B1(n801), .B2(n1548), .A(n1547), .ZN(n1637) );
  INV_X1 U1698 ( .A(n1637), .ZN(n1676) );
  NOR2_X1 U1699 ( .A1(n806), .A2(n1676), .ZN(normResult[2]) );
  OAI22_X1 U1700 ( .A1(n23), .A2(n1549), .B1(n1678), .B2(n1548), .ZN(n1673) );
  INV_X1 U1701 ( .A(n1673), .ZN(n1639) );
  OAI22_X1 U1702 ( .A1(n268), .A2(n1552), .B1(n1551), .B2(n1550), .ZN(n1664)
         );
  INV_X1 U1703 ( .A(n1664), .ZN(n1588) );
  OAI22_X1 U1704 ( .A1(n147), .A2(n1556), .B1(n1555), .B2(n1554), .ZN(n1655)
         );
  INV_X1 U1705 ( .A(n1655), .ZN(n1578) );
  INV_X1 U1706 ( .A(n1682), .ZN(n1559) );
  OAI22_X1 U1707 ( .A1(n85), .A2(n1560), .B1(n1559), .B2(n379), .ZN(n1645) );
  INV_X1 U1708 ( .A(n1645), .ZN(n1568) );
  INV_X1 U1709 ( .A(n1616), .ZN(n1686) );
  INV_X1 U1710 ( .A(n223), .ZN(n1646) );
  AOI22_X1 U1711 ( .A1(n1646), .A2(n1565), .B1(n1564), .B2(n1563), .ZN(n1566)
         );
  OAI221_X1 U1712 ( .B1(n158), .B2(n1568), .C1(n1686), .C2(n1567), .A(n1566), 
        .ZN(n1570) );
  INV_X1 U1713 ( .A(n1570), .ZN(n1691) );
  OAI222_X1 U1714 ( .A1(n1653), .A2(n814), .B1(n811), .B2(n1691), .C1(n246), 
        .C2(n1571), .ZN(n1725) );
  INV_X1 U1715 ( .A(n1725), .ZN(n1694) );
  INV_X1 U1716 ( .A(n619), .ZN(n1656) );
  AOI22_X1 U1717 ( .A1(n1656), .A2(n1575), .B1(n558), .B2(n1573), .ZN(n1576)
         );
  OAI221_X1 U1718 ( .B1(n1579), .B2(n1578), .C1(n1694), .C2(n1577), .A(n1576), 
        .ZN(n1580) );
  INV_X1 U1719 ( .A(n1580), .ZN(n1696) );
  OAI222_X1 U1720 ( .A1(n1662), .A2(n815), .B1(n823), .B2(n1696), .C1(n397), 
        .C2(n1581), .ZN(n1730) );
  INV_X1 U1721 ( .A(n1730), .ZN(n1699) );
  INV_X1 U1722 ( .A(n475), .ZN(n1665) );
  AOI22_X1 U1723 ( .A1(n1665), .A2(n1585), .B1(n749), .B2(n1583), .ZN(n1586)
         );
  OAI221_X1 U1724 ( .B1(n252), .B2(n1588), .C1(n1699), .C2(n1587), .A(n1586), 
        .ZN(n1590) );
  INV_X1 U1725 ( .A(n1590), .ZN(n1701) );
  OAI222_X1 U1726 ( .A1(n1671), .A2(n816), .B1(n824), .B2(n1701), .C1(n366), 
        .C2(n1591), .ZN(n1735) );
  INV_X1 U1727 ( .A(n1735), .ZN(n1704) );
  NAND2_X1 U1728 ( .A1(n478), .A2(n642), .ZN(n1643) );
  INV_X1 U1729 ( .A(n1596), .ZN(n1593) );
  OAI21_X1 U1730 ( .B1(n559), .B2(n1593), .A(n43), .ZN(n1595) );
  INV_X1 U1731 ( .A(n1595), .ZN(n1902) );
  OAI21_X1 U1732 ( .B1(n1597), .B2(n1641), .A(n35), .ZN(n1598) );
  INV_X1 U1733 ( .A(n34), .ZN(n1899) );
  INV_X1 U1734 ( .A(n103), .ZN(n1603) );
  NAND2_X1 U1735 ( .A1(n539), .A2(n480), .ZN(n1610) );
  INV_X1 U1736 ( .A(n1610), .ZN(n1607) );
  INV_X1 U1737 ( .A(n329), .ZN(n1602) );
  OAI21_X1 U1738 ( .B1(n709), .B2(n45), .A(n1604), .ZN(n1605) );
  INV_X1 U1739 ( .A(n1605), .ZN(n1913) );
  OAI21_X1 U1740 ( .B1(n1607), .B2(n56), .A(n1606), .ZN(n1609) );
  INV_X1 U1741 ( .A(n1609), .ZN(n1910) );
  OAI21_X1 U1742 ( .B1(n480), .B2(n317), .A(n1610), .ZN(n1612) );
  INV_X1 U1743 ( .A(n1612), .ZN(n1907) );
  INV_X1 U1744 ( .A(n481), .ZN(n1905) );
  INV_X1 U1745 ( .A(n1839), .ZN(n1855) );
  INV_X1 U1746 ( .A(n1765), .ZN(n1787) );
  INV_X1 U1747 ( .A(n1648), .ZN(n1688) );
  AOI222_X1 U1748 ( .A1(n1616), .A2(n695), .B1(n198), .B2(n1684), .C1(n1681), 
        .C2(n1615), .ZN(n1617) );
  OAI221_X1 U1749 ( .B1(n1689), .B2(n1618), .C1(n1687), .C2(n1688), .A(n1617), 
        .ZN(n1619) );
  INV_X1 U1750 ( .A(n1619), .ZN(n1724) );
  OAI222_X1 U1751 ( .A1(n1719), .A2(n814), .B1(n1724), .B2(n246), .C1(n812), 
        .C2(n1620), .ZN(n1783) );
  AOI222_X1 U1752 ( .A1(n1764), .A2(n631), .B1(n641), .B2(n1783), .C1(n1780), 
        .C2(n1621), .ZN(n1622) );
  OAI221_X1 U1753 ( .B1(n1788), .B2(n1623), .C1(n1786), .C2(n1787), .A(n1622), 
        .ZN(n1624) );
  INV_X1 U1754 ( .A(n1624), .ZN(n1813) );
  OAI222_X1 U1755 ( .A1(n1808), .A2(n815), .B1(n1813), .B2(n397), .C1(n823), 
        .C2(n1625), .ZN(n1851) );
  AOI222_X1 U1756 ( .A1(n1838), .A2(n730), .B1(n315), .B2(n1851), .C1(n1849), 
        .C2(n1626), .ZN(n1627) );
  OAI221_X1 U1757 ( .B1(n1856), .B2(n1628), .C1(n1854), .C2(n1855), .A(n1627), 
        .ZN(n1629) );
  INV_X1 U1758 ( .A(n1629), .ZN(n1871) );
  OAI222_X1 U1759 ( .A1(n1866), .A2(n816), .B1(n1871), .B2(n366), .C1(n824), 
        .C2(n1630), .ZN(n1891) );
  OAI22_X1 U1760 ( .A1(n1678), .A2(n1889), .B1(n802), .B2(n1631), .ZN(n1890)
         );
  NAND2_X1 U1761 ( .A1(n63), .A2(n806), .ZN(n1896) );
  INV_X1 U1762 ( .A(n474), .ZN(n1898) );
  INV_X1 U1763 ( .A(n1635), .ZN(n1636) );
  AOI22_X1 U1764 ( .A1(n442), .A2(n1637), .B1(n748), .B2(n1636), .ZN(n1638) );
  OAI221_X1 U1765 ( .B1(n806), .B2(n1639), .C1(n1704), .C2(n1643), .A(n1638), 
        .ZN(normResult[3]) );
  OAI22_X1 U1766 ( .A1(n1678), .A2(n806), .B1(n802), .B2(n1896), .ZN(n1642) );
  INV_X1 U1767 ( .A(n1644), .ZN(n1647) );
  AOI222_X1 U1768 ( .A1(n1681), .A2(n1648), .B1(n1647), .B2(n1684), .C1(n1646), 
        .C2(n1645), .ZN(n1649) );
  OAI221_X1 U1769 ( .B1(n1689), .B2(n1686), .C1(n1651), .C2(n541), .A(n1649), 
        .ZN(n1652) );
  INV_X1 U1770 ( .A(n1652), .ZN(n1705) );
  OAI222_X1 U1771 ( .A1(n1691), .A2(n814), .B1(n812), .B2(n1705), .C1(n1653), 
        .C2(n246), .ZN(n1738) );
  INV_X1 U1772 ( .A(n1654), .ZN(n1657) );
  AOI222_X1 U1773 ( .A1(n1780), .A2(n1738), .B1(n1657), .B2(n1706), .C1(n1656), 
        .C2(n1655), .ZN(n1658) );
  OAI221_X1 U1774 ( .B1(n1788), .B2(n1694), .C1(n1660), .C2(n620), .A(n1658), 
        .ZN(n1661) );
  INV_X1 U1775 ( .A(n1661), .ZN(n1710) );
  OAI222_X1 U1776 ( .A1(n1696), .A2(n815), .B1(n823), .B2(n1710), .C1(n1662), 
        .C2(n397), .ZN(n1743) );
  INV_X1 U1777 ( .A(n1663), .ZN(n1666) );
  AOI222_X1 U1778 ( .A1(n1849), .A2(n1743), .B1(n1666), .B2(n1711), .C1(n1665), 
        .C2(n1664), .ZN(n1667) );
  OAI221_X1 U1779 ( .B1(n1856), .B2(n1699), .C1(n1669), .C2(n378), .A(n1667), 
        .ZN(n1670) );
  INV_X1 U1780 ( .A(n1670), .ZN(n1715) );
  OAI222_X1 U1781 ( .A1(n1701), .A2(n817), .B1(n824), .B2(n1715), .C1(n1671), 
        .C2(n366), .ZN(n1748) );
  INV_X1 U1782 ( .A(n1886), .ZN(n1674) );
  AOI222_X1 U1783 ( .A1(n1883), .A2(n1748), .B1(n1674), .B2(n1716), .C1(n442), 
        .C2(n1673), .ZN(n1675) );
  OAI221_X1 U1784 ( .B1(n1888), .B2(n1704), .C1(n1676), .C2(n520), .A(n1675), 
        .ZN(normResult[4]) );
  INV_X1 U1785 ( .A(n1748), .ZN(n1718) );
  INV_X1 U1786 ( .A(n1743), .ZN(n1713) );
  INV_X1 U1787 ( .A(n1738), .ZN(n1708) );
  AOI222_X1 U1788 ( .A1(n1684), .A2(n695), .B1(n198), .B2(n1682), .C1(n1681), 
        .C2(n1680), .ZN(n1685) );
  OAI221_X1 U1789 ( .B1(n1689), .B2(n1688), .C1(n1687), .C2(n1686), .A(n1685), 
        .ZN(n1690) );
  INV_X1 U1790 ( .A(n1690), .ZN(n1722) );
  OAI222_X1 U1791 ( .A1(n1705), .A2(n814), .B1(n812), .B2(n1722), .C1(n1691), 
        .C2(n246), .ZN(n1751) );
  AOI222_X1 U1792 ( .A1(n1706), .A2(n679), .B1(n1692), .B2(n641), .C1(n1780), 
        .C2(n1751), .ZN(n1693) );
  OAI221_X1 U1793 ( .B1(n1788), .B2(n1708), .C1(n1786), .C2(n1694), .A(n1693), 
        .ZN(n1695) );
  INV_X1 U1794 ( .A(n1695), .ZN(n1729) );
  OAI222_X1 U1795 ( .A1(n1710), .A2(n815), .B1(n823), .B2(n1729), .C1(n1696), 
        .C2(n397), .ZN(n1756) );
  AOI222_X1 U1796 ( .A1(n1711), .A2(n730), .B1(n1697), .B2(n315), .C1(n1849), 
        .C2(n1756), .ZN(n1698) );
  OAI221_X1 U1797 ( .B1(n1856), .B2(n1713), .C1(n1854), .C2(n1699), .A(n1698), 
        .ZN(n1700) );
  INV_X1 U1798 ( .A(n1700), .ZN(n1734) );
  OAI222_X1 U1799 ( .A1(n1715), .A2(n817), .B1(n824), .B2(n1734), .C1(n1701), 
        .C2(n366), .ZN(n1761) );
  AOI222_X1 U1800 ( .A1(n1716), .A2(n64), .B1(n1702), .B2(n94), .C1(n1883), 
        .C2(n1761), .ZN(n1703) );
  INV_X1 U1801 ( .A(n1761), .ZN(n1737) );
  INV_X1 U1802 ( .A(n1756), .ZN(n1732) );
  INV_X1 U1803 ( .A(n1751), .ZN(n1727) );
  AOI222_X1 U1804 ( .A1(n1725), .A2(n631), .B1(n641), .B2(n1706), .C1(n1780), 
        .C2(n1766), .ZN(n1707) );
  OAI221_X1 U1805 ( .B1(n1788), .B2(n1727), .C1(n1786), .C2(n1708), .A(n1707), 
        .ZN(n1709) );
  INV_X1 U1806 ( .A(n1709), .ZN(n1742) );
  OAI222_X1 U1807 ( .A1(n1729), .A2(n815), .B1(n823), .B2(n1742), .C1(n1710), 
        .C2(n397), .ZN(n1771) );
  AOI222_X1 U1808 ( .A1(n1730), .A2(n730), .B1(n315), .B2(n1711), .C1(n1849), 
        .C2(n1771), .ZN(n1712) );
  OAI221_X1 U1809 ( .B1(n1856), .B2(n1732), .C1(n1854), .C2(n1713), .A(n1712), 
        .ZN(n1714) );
  INV_X1 U1810 ( .A(n1714), .ZN(n1747) );
  AOI222_X1 U1811 ( .A1(n1892), .A2(n1735), .B1(n94), .B2(n1716), .C1(n1883), 
        .C2(n1776), .ZN(n1717) );
  OAI221_X1 U1812 ( .B1(n1888), .B2(n1737), .C1(n1718), .C2(n1886), .A(n1717), 
        .ZN(normResult[6]) );
  INV_X1 U1813 ( .A(n1776), .ZN(n1750) );
  INV_X1 U1814 ( .A(n1771), .ZN(n1745) );
  INV_X1 U1815 ( .A(n1766), .ZN(n1740) );
  OAI222_X1 U1816 ( .A1(n1724), .A2(n814), .B1(n1722), .B2(n246), .C1(n812), 
        .C2(n1719), .ZN(n1781) );
  AOI222_X1 U1817 ( .A1(n1738), .A2(n679), .B1(n641), .B2(n1725), .C1(n1780), 
        .C2(n1781), .ZN(n1726) );
  OAI221_X1 U1818 ( .B1(n1788), .B2(n1740), .C1(n1786), .C2(n1727), .A(n1726), 
        .ZN(n1728) );
  INV_X1 U1819 ( .A(n1728), .ZN(n1755) );
  OAI222_X1 U1820 ( .A1(n1742), .A2(n815), .B1(n823), .B2(n1755), .C1(n1729), 
        .C2(n397), .ZN(n1791) );
  AOI222_X1 U1821 ( .A1(n1743), .A2(n730), .B1(n315), .B2(n1730), .C1(n1849), 
        .C2(n1791), .ZN(n1731) );
  OAI221_X1 U1822 ( .B1(n1856), .B2(n1745), .C1(n1854), .C2(n1732), .A(n1731), 
        .ZN(n1733) );
  INV_X1 U1823 ( .A(n1733), .ZN(n1760) );
  AOI222_X1 U1824 ( .A1(n1748), .A2(n64), .B1(n94), .B2(n1735), .C1(n1883), 
        .C2(n1796), .ZN(n1736) );
  INV_X1 U1825 ( .A(n1796), .ZN(n1763) );
  INV_X1 U1826 ( .A(n1791), .ZN(n1758) );
  INV_X1 U1827 ( .A(n1781), .ZN(n1753) );
  AOI222_X1 U1828 ( .A1(n1751), .A2(n631), .B1(n641), .B2(n1738), .C1(n1780), 
        .C2(n1783), .ZN(n1739) );
  OAI221_X1 U1829 ( .B1(n1788), .B2(n1753), .C1(n1786), .C2(n1740), .A(n1739), 
        .ZN(n1741) );
  INV_X1 U1830 ( .A(n1741), .ZN(n1770) );
  OAI222_X1 U1831 ( .A1(n1755), .A2(n815), .B1(n823), .B2(n1770), .C1(n1742), 
        .C2(n397), .ZN(n1800) );
  AOI222_X1 U1832 ( .A1(n1756), .A2(n730), .B1(n315), .B2(n1743), .C1(n1849), 
        .C2(n1800), .ZN(n1744) );
  OAI221_X1 U1833 ( .B1(n1856), .B2(n1758), .C1(n1854), .C2(n1745), .A(n1744), 
        .ZN(n1746) );
  INV_X1 U1834 ( .A(n1746), .ZN(n1775) );
  OAI222_X1 U1835 ( .A1(n1760), .A2(n817), .B1(n824), .B2(n1775), .C1(n1747), 
        .C2(n366), .ZN(n1805) );
  AOI222_X1 U1836 ( .A1(n1761), .A2(n1892), .B1(n94), .B2(n1748), .C1(n1883), 
        .C2(n1805), .ZN(n1749) );
  INV_X1 U1837 ( .A(n1805), .ZN(n1778) );
  INV_X1 U1838 ( .A(n1800), .ZN(n1773) );
  INV_X1 U1839 ( .A(n1783), .ZN(n1768) );
  AOI222_X1 U1840 ( .A1(n1766), .A2(n679), .B1(n641), .B2(n1751), .C1(n1780), 
        .C2(n1764), .ZN(n1752) );
  OAI221_X1 U1841 ( .B1(n1788), .B2(n1768), .C1(n1786), .C2(n1753), .A(n1752), 
        .ZN(n1754) );
  INV_X1 U1842 ( .A(n1754), .ZN(n1790) );
  OAI222_X1 U1843 ( .A1(n1770), .A2(n815), .B1(n823), .B2(n1790), .C1(n1755), 
        .C2(n397), .ZN(n1814) );
  AOI222_X1 U1844 ( .A1(n1771), .A2(n730), .B1(n315), .B2(n1756), .C1(n1849), 
        .C2(n1814), .ZN(n1757) );
  OAI221_X1 U1845 ( .B1(n1856), .B2(n1773), .C1(n1854), .C2(n1758), .A(n1757), 
        .ZN(n1759) );
  INV_X1 U1846 ( .A(n1759), .ZN(n1795) );
  OAI222_X1 U1847 ( .A1(n1775), .A2(n817), .B1(n824), .B2(n1795), .C1(n1760), 
        .C2(n366), .ZN(n1819) );
  AOI222_X1 U1848 ( .A1(n1776), .A2(n64), .B1(n94), .B2(n1761), .C1(n1883), 
        .C2(n1819), .ZN(n1762) );
  OAI221_X1 U1849 ( .B1(n1888), .B2(n1778), .C1(n1763), .C2(n1886), .A(n1762), 
        .ZN(normResult[9]) );
  INV_X1 U1850 ( .A(n1819), .ZN(n1798) );
  INV_X1 U1851 ( .A(n1814), .ZN(n1793) );
  INV_X1 U1852 ( .A(n1764), .ZN(n1785) );
  AOI222_X1 U1853 ( .A1(n1781), .A2(n631), .B1(n641), .B2(n1766), .C1(n1780), 
        .C2(n1765), .ZN(n1767) );
  OAI221_X1 U1854 ( .B1(n1788), .B2(n1785), .C1(n1786), .C2(n1768), .A(n1767), 
        .ZN(n1769) );
  INV_X1 U1855 ( .A(n1769), .ZN(n1799) );
  OAI222_X1 U1856 ( .A1(n1790), .A2(n815), .B1(n823), .B2(n1799), .C1(n1770), 
        .C2(n397), .ZN(n1822) );
  AOI222_X1 U1857 ( .A1(n1791), .A2(n730), .B1(n315), .B2(n1771), .C1(n1849), 
        .C2(n1822), .ZN(n1772) );
  OAI221_X1 U1858 ( .B1(n1856), .B2(n1793), .C1(n1854), .C2(n1773), .A(n1772), 
        .ZN(n1774) );
  INV_X1 U1859 ( .A(n1774), .ZN(n1804) );
  OAI222_X1 U1860 ( .A1(n1795), .A2(n816), .B1(n824), .B2(n1804), .C1(n1775), 
        .C2(n366), .ZN(n1827) );
  AOI222_X1 U1861 ( .A1(n1796), .A2(n1892), .B1(n94), .B2(n1776), .C1(n1883), 
        .C2(n1827), .ZN(n1777) );
  INV_X1 U1862 ( .A(n1827), .ZN(n1807) );
  INV_X1 U1863 ( .A(n1822), .ZN(n1802) );
  AOI222_X1 U1864 ( .A1(n1783), .A2(n679), .B1(n641), .B2(n1781), .C1(n1780), 
        .C2(n1779), .ZN(n1784) );
  OAI221_X1 U1865 ( .B1(n1788), .B2(n1787), .C1(n1786), .C2(n1785), .A(n1784), 
        .ZN(n1789) );
  INV_X1 U1866 ( .A(n1789), .ZN(n1811) );
  OAI222_X1 U1867 ( .A1(n1799), .A2(n815), .B1(n823), .B2(n1811), .C1(n1790), 
        .C2(n397), .ZN(n1830) );
  AOI222_X1 U1868 ( .A1(n1800), .A2(n730), .B1(n315), .B2(n1791), .C1(n1849), 
        .C2(n1830), .ZN(n1792) );
  OAI221_X1 U1869 ( .B1(n1856), .B2(n1802), .C1(n1854), .C2(n1793), .A(n1792), 
        .ZN(n1794) );
  INV_X1 U1870 ( .A(n1794), .ZN(n1818) );
  OAI222_X1 U1871 ( .A1(n1804), .A2(n816), .B1(n824), .B2(n1818), .C1(n1795), 
        .C2(n366), .ZN(n1835) );
  AOI222_X1 U1872 ( .A1(n1805), .A2(n1892), .B1(n94), .B2(n1796), .C1(n1883), 
        .C2(n1835), .ZN(n1797) );
  OAI221_X1 U1873 ( .B1(n1888), .B2(n1807), .C1(n1798), .C2(n1886), .A(n1797), 
        .ZN(normResult[11]) );
  INV_X1 U1874 ( .A(n1835), .ZN(n1821) );
  INV_X1 U1875 ( .A(n1830), .ZN(n1816) );
  AOI222_X1 U1876 ( .A1(n1814), .A2(n730), .B1(n315), .B2(n1800), .C1(n1849), 
        .C2(n1840), .ZN(n1801) );
  OAI221_X1 U1877 ( .B1(n1856), .B2(n1816), .C1(n1854), .C2(n1802), .A(n1801), 
        .ZN(n1803) );
  INV_X1 U1878 ( .A(n1803), .ZN(n1826) );
  OAI222_X1 U1879 ( .A1(n1818), .A2(n817), .B1(n824), .B2(n1826), .C1(n1804), 
        .C2(n366), .ZN(n1845) );
  AOI222_X1 U1880 ( .A1(n1819), .A2(n1892), .B1(n791), .B2(n1805), .C1(n1883), 
        .C2(n1845), .ZN(n1806) );
  OAI221_X1 U1881 ( .B1(n1888), .B2(n1821), .C1(n1807), .C2(n1886), .A(n1806), 
        .ZN(normResult[12]) );
  INV_X1 U1882 ( .A(n1845), .ZN(n1829) );
  INV_X1 U1883 ( .A(n1840), .ZN(n1824) );
  OAI222_X1 U1884 ( .A1(n1813), .A2(n815), .B1(n1811), .B2(n397), .C1(n823), 
        .C2(n1808), .ZN(n1850) );
  AOI222_X1 U1885 ( .A1(n1822), .A2(n730), .B1(n315), .B2(n1814), .C1(n1849), 
        .C2(n1850), .ZN(n1815) );
  OAI221_X1 U1886 ( .B1(n1856), .B2(n1824), .C1(n1854), .C2(n1816), .A(n1815), 
        .ZN(n1817) );
  INV_X1 U1887 ( .A(n1817), .ZN(n1834) );
  OAI222_X1 U1888 ( .A1(n1826), .A2(n817), .B1(n824), .B2(n1834), .C1(n1818), 
        .C2(n366), .ZN(n1859) );
  AOI222_X1 U1889 ( .A1(n1827), .A2(n64), .B1(n791), .B2(n1819), .C1(n1883), 
        .C2(n1859), .ZN(n1820) );
  OAI221_X1 U1890 ( .B1(n1888), .B2(n1829), .C1(n1821), .C2(n1886), .A(n1820), 
        .ZN(normResult[13]) );
  INV_X1 U1891 ( .A(n1859), .ZN(n1837) );
  INV_X1 U1892 ( .A(n1850), .ZN(n1832) );
  AOI222_X1 U1893 ( .A1(n1830), .A2(n730), .B1(n315), .B2(n1822), .C1(n1849), 
        .C2(n1851), .ZN(n1823) );
  OAI221_X1 U1894 ( .B1(n1856), .B2(n1832), .C1(n1854), .C2(n1824), .A(n1823), 
        .ZN(n1825) );
  INV_X1 U1895 ( .A(n1825), .ZN(n1844) );
  OAI222_X1 U1896 ( .A1(n1834), .A2(n816), .B1(n824), .B2(n1844), .C1(n1826), 
        .C2(n366), .ZN(n1863) );
  AOI222_X1 U1897 ( .A1(n1835), .A2(n64), .B1(n791), .B2(n1827), .C1(n1883), 
        .C2(n1863), .ZN(n1828) );
  OAI221_X1 U1898 ( .B1(n1888), .B2(n1837), .C1(n1829), .C2(n1886), .A(n1828), 
        .ZN(normResult[14]) );
  INV_X1 U1899 ( .A(n1863), .ZN(n1847) );
  INV_X1 U1900 ( .A(n1851), .ZN(n1842) );
  AOI222_X1 U1901 ( .A1(n1840), .A2(n730), .B1(n315), .B2(n1830), .C1(n1849), 
        .C2(n1838), .ZN(n1831) );
  OAI221_X1 U1902 ( .B1(n1856), .B2(n1842), .C1(n1854), .C2(n1832), .A(n1831), 
        .ZN(n1833) );
  INV_X1 U1903 ( .A(n1833), .ZN(n1858) );
  OAI222_X1 U1904 ( .A1(n1844), .A2(n816), .B1(n824), .B2(n1858), .C1(n1834), 
        .C2(n366), .ZN(n1872) );
  AOI222_X1 U1905 ( .A1(n1845), .A2(n1892), .B1(n791), .B2(n1835), .C1(n1883), 
        .C2(n1872), .ZN(n1836) );
  OAI221_X1 U1906 ( .B1(n1888), .B2(n1847), .C1(n1837), .C2(n1886), .A(n1836), 
        .ZN(normResult[15]) );
  INV_X1 U1907 ( .A(n1872), .ZN(n1861) );
  INV_X1 U1908 ( .A(n1838), .ZN(n1853) );
  AOI222_X1 U1909 ( .A1(n1850), .A2(n730), .B1(n315), .B2(n1840), .C1(n1849), 
        .C2(n1839), .ZN(n1841) );
  OAI221_X1 U1910 ( .B1(n1856), .B2(n1853), .C1(n1854), .C2(n1842), .A(n1841), 
        .ZN(n1843) );
  INV_X1 U1911 ( .A(n1843), .ZN(n1862) );
  OAI222_X1 U1912 ( .A1(n1858), .A2(n817), .B1(n824), .B2(n1862), .C1(n1844), 
        .C2(n366), .ZN(n1875) );
  AOI222_X1 U1913 ( .A1(n1859), .A2(n1892), .B1(n791), .B2(n1845), .C1(n1883), 
        .C2(n1875), .ZN(n1846) );
  OAI221_X1 U1914 ( .B1(n1888), .B2(n1861), .C1(n1847), .C2(n1886), .A(n1846), 
        .ZN(normResult[16]) );
  INV_X1 U1915 ( .A(n1875), .ZN(n1865) );
  AOI222_X1 U1916 ( .A1(n1851), .A2(n730), .B1(n315), .B2(n1850), .C1(n1849), 
        .C2(n1848), .ZN(n1852) );
  OAI221_X1 U1917 ( .B1(n1856), .B2(n1855), .C1(n1854), .C2(n1853), .A(n1852), 
        .ZN(n1857) );
  INV_X1 U1918 ( .A(n1857), .ZN(n1869) );
  OAI222_X1 U1919 ( .A1(n1862), .A2(n817), .B1(n824), .B2(n1869), .C1(n1858), 
        .C2(n366), .ZN(n1879) );
  AOI222_X1 U1920 ( .A1(n1863), .A2(n64), .B1(n791), .B2(n1859), .C1(n1883), 
        .C2(n1879), .ZN(n1860) );
  OAI221_X1 U1921 ( .B1(n1888), .B2(n1865), .C1(n1861), .C2(n1886), .A(n1860), 
        .ZN(normResult[17]) );
  INV_X1 U1922 ( .A(n1879), .ZN(n1874) );
  OAI222_X1 U1923 ( .A1(n1862), .A2(n366), .B1(n1869), .B2(n817), .C1(n824), 
        .C2(n1871), .ZN(n1884) );
  AOI222_X1 U1924 ( .A1(n1872), .A2(n64), .B1(n791), .B2(n1863), .C1(n1883), 
        .C2(n1884), .ZN(n1864) );
  OAI221_X1 U1925 ( .B1(n1888), .B2(n1874), .C1(n1865), .C2(n1886), .A(n1864), 
        .ZN(normResult[18]) );
  INV_X1 U1926 ( .A(n1884), .ZN(n1877) );
  AOI222_X1 U1927 ( .A1(n1875), .A2(n64), .B1(n791), .B2(n1872), .C1(n1883), 
        .C2(n1893), .ZN(n1873) );
  OAI221_X1 U1928 ( .B1(n1877), .B2(n1888), .C1(n1874), .C2(n1886), .A(n1873), 
        .ZN(normResult[19]) );
  INV_X1 U1929 ( .A(n1893), .ZN(n1881) );
  AOI222_X1 U1930 ( .A1(n1879), .A2(n64), .B1(n791), .B2(n1875), .C1(n1883), 
        .C2(n1891), .ZN(n1876) );
  OAI221_X1 U1931 ( .B1(n1881), .B2(n1888), .C1(n1877), .C2(n1886), .A(n1876), 
        .ZN(normResult[20]) );
  INV_X1 U1932 ( .A(n1891), .ZN(n1887) );
  AOI222_X1 U1933 ( .A1(n1884), .A2(n64), .B1(n791), .B2(n1879), .C1(n1883), 
        .C2(n1878), .ZN(n1880) );
  OAI221_X1 U1934 ( .B1(n1887), .B2(n1888), .C1(n1881), .C2(n1886), .A(n1880), 
        .ZN(normResult[21]) );
  AOI222_X1 U1935 ( .A1(n1892), .A2(n1893), .B1(n791), .B2(n1884), .C1(n1883), 
        .C2(n1882), .ZN(n1885) );
  OAI221_X1 U1936 ( .B1(n1889), .B2(n1888), .C1(n1887), .C2(n1886), .A(n1885), 
        .ZN(normResult[22]) );
  INV_X1 U1937 ( .A(n1890), .ZN(n1897) );
  AOI22_X1 U1938 ( .A1(n94), .A2(n1893), .B1(n64), .B2(n1891), .ZN(n1894) );
  OAI211_X1 U1939 ( .C1(n1897), .C2(n462), .A(n1895), .B(n1894), .ZN(
        normResult[23]) );
  OAI21_X1 U1940 ( .B1(n1899), .B2(n748), .A(n1900), .ZN(normExponent[0]) );
  INV_X1 U1941 ( .A(n1900), .ZN(n1901) );
  OAI21_X1 U1942 ( .B1(n1902), .B2(n1901), .A(n1903), .ZN(normExponent[1]) );
  INV_X1 U1943 ( .A(n1903), .ZN(n1904) );
  OAI21_X1 U1944 ( .B1(n1904), .B2(n1905), .A(n1906), .ZN(normExponent[2]) );
  NAND2_X1 U1945 ( .A1(n594), .A2(n1907), .ZN(n1908) );
  OAI21_X1 U1946 ( .B1(n1907), .B2(n594), .A(n1908), .ZN(normExponent[3]) );
  INV_X1 U1947 ( .A(n1908), .ZN(n1909) );
  OAI21_X1 U1948 ( .B1(n40), .B2(n1909), .A(n384), .ZN(normExponent[4]) );
  INV_X1 U1949 ( .A(n384), .ZN(n1912) );
  OAI21_X1 U1950 ( .B1(n479), .B2(n1912), .A(n352), .ZN(normExponent[5]) );
  INV_X1 U1951 ( .A(n352), .ZN(n1917) );
  AOI21_X1 U1952 ( .B1(n1917), .B2(n647), .A(n25), .ZN(normExponent[7]) );
endmodule


module FPAdder ( clk, a, b, result, overflow, underflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input clk;
  output overflow, underflow;
  wire   f_bigger, signFO, signSO, finalSign, cout, N30, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4;
  wire   [31:23] a_reg;
  wire   [22:0] a_whole;
  wire   [31:23] b_reg;
  wire   [22:0] b_whole;
  wire   [4:0] shiftAmount;
  wire   [23:0] shiftedResult;
  wire   [23:0] tempResult;
  wire   [7:0] outputExponent;
  wire   [22:0] normResult;

  DFF_X1 a_reg_reg_31_ ( .D(a[31]), .CK(clk), .Q(a_reg[31]) );
  DFF_X1 a_reg_reg_30_ ( .D(a[30]), .CK(clk), .Q(a_reg[30]) );
  DFF_X1 a_reg_reg_29_ ( .D(a[29]), .CK(clk), .Q(a_reg[29]) );
  DFF_X1 a_reg_reg_28_ ( .D(a[28]), .CK(clk), .Q(a_reg[28]) );
  DFF_X1 a_reg_reg_27_ ( .D(a[27]), .CK(clk), .Q(a_reg[27]) );
  DFF_X1 a_reg_reg_26_ ( .D(a[26]), .CK(clk), .Q(a_reg[26]) );
  DFF_X1 a_reg_reg_25_ ( .D(a[25]), .CK(clk), .Q(a_reg[25]) );
  DFF_X1 a_reg_reg_24_ ( .D(a[24]), .CK(clk), .Q(a_reg[24]) );
  DFF_X1 a_reg_reg_23_ ( .D(a[23]), .CK(clk), .Q(a_reg[23]) );
  DFF_X1 a_reg_reg_22_ ( .D(a[22]), .CK(clk), .Q(a_whole[22]) );
  DFF_X1 a_reg_reg_21_ ( .D(a[21]), .CK(clk), .Q(a_whole[21]) );
  DFF_X1 a_reg_reg_20_ ( .D(a[20]), .CK(clk), .Q(a_whole[20]) );
  DFF_X1 a_reg_reg_19_ ( .D(a[19]), .CK(clk), .Q(a_whole[19]) );
  DFF_X1 a_reg_reg_18_ ( .D(a[18]), .CK(clk), .Q(a_whole[18]) );
  DFF_X1 a_reg_reg_17_ ( .D(a[17]), .CK(clk), .Q(a_whole[17]) );
  DFF_X1 a_reg_reg_16_ ( .D(a[16]), .CK(clk), .Q(a_whole[16]) );
  DFF_X1 a_reg_reg_15_ ( .D(a[15]), .CK(clk), .Q(a_whole[15]) );
  DFF_X1 a_reg_reg_14_ ( .D(a[14]), .CK(clk), .Q(a_whole[14]) );
  DFF_X1 a_reg_reg_13_ ( .D(a[13]), .CK(clk), .Q(a_whole[13]) );
  DFF_X1 a_reg_reg_12_ ( .D(a[12]), .CK(clk), .Q(a_whole[12]) );
  DFF_X1 a_reg_reg_11_ ( .D(a[11]), .CK(clk), .Q(a_whole[11]) );
  DFF_X1 a_reg_reg_10_ ( .D(a[10]), .CK(clk), .Q(a_whole[10]) );
  DFF_X1 a_reg_reg_9_ ( .D(a[9]), .CK(clk), .Q(a_whole[9]) );
  DFF_X1 a_reg_reg_8_ ( .D(a[8]), .CK(clk), .Q(a_whole[8]) );
  DFF_X1 a_reg_reg_7_ ( .D(a[7]), .CK(clk), .Q(a_whole[7]) );
  DFF_X1 a_reg_reg_6_ ( .D(a[6]), .CK(clk), .Q(a_whole[6]) );
  DFF_X1 a_reg_reg_5_ ( .D(a[5]), .CK(clk), .Q(a_whole[5]) );
  DFF_X1 a_reg_reg_4_ ( .D(a[4]), .CK(clk), .Q(a_whole[4]) );
  DFF_X1 a_reg_reg_3_ ( .D(a[3]), .CK(clk), .Q(a_whole[3]) );
  DFF_X1 a_reg_reg_2_ ( .D(a[2]), .CK(clk), .Q(a_whole[2]) );
  DFF_X1 a_reg_reg_1_ ( .D(a[1]), .CK(clk), .Q(a_whole[1]) );
  DFF_X1 a_reg_reg_0_ ( .D(a[0]), .CK(clk), .Q(a_whole[0]) );
  DFF_X1 b_reg_reg_31_ ( .D(b[31]), .CK(clk), .Q(b_reg[31]) );
  DFF_X1 b_reg_reg_30_ ( .D(b[30]), .CK(clk), .Q(b_reg[30]) );
  DFF_X1 b_reg_reg_29_ ( .D(b[29]), .CK(clk), .Q(b_reg[29]) );
  DFF_X1 b_reg_reg_28_ ( .D(b[28]), .CK(clk), .Q(b_reg[28]) );
  DFF_X1 b_reg_reg_27_ ( .D(b[27]), .CK(clk), .Q(b_reg[27]) );
  DFF_X1 b_reg_reg_26_ ( .D(b[26]), .CK(clk), .Q(b_reg[26]) );
  DFF_X1 b_reg_reg_25_ ( .D(b[25]), .CK(clk), .Q(b_reg[25]) );
  DFF_X1 b_reg_reg_24_ ( .D(b[24]), .CK(clk), .Q(b_reg[24]) );
  DFF_X1 b_reg_reg_23_ ( .D(b[23]), .CK(clk), .Q(b_reg[23]) );
  DFF_X1 b_reg_reg_22_ ( .D(b[22]), .CK(clk), .Q(b_whole[22]) );
  DFF_X1 b_reg_reg_21_ ( .D(b[21]), .CK(clk), .Q(b_whole[21]) );
  DFF_X1 b_reg_reg_20_ ( .D(b[20]), .CK(clk), .Q(b_whole[20]) );
  DFF_X1 b_reg_reg_19_ ( .D(b[19]), .CK(clk), .Q(b_whole[19]) );
  DFF_X1 b_reg_reg_18_ ( .D(b[18]), .CK(clk), .Q(b_whole[18]) );
  DFF_X1 b_reg_reg_17_ ( .D(b[17]), .CK(clk), .Q(b_whole[17]) );
  DFF_X1 b_reg_reg_16_ ( .D(b[16]), .CK(clk), .Q(b_whole[16]) );
  DFF_X1 b_reg_reg_15_ ( .D(b[15]), .CK(clk), .Q(b_whole[15]) );
  DFF_X1 b_reg_reg_14_ ( .D(b[14]), .CK(clk), .Q(b_whole[14]) );
  DFF_X1 b_reg_reg_13_ ( .D(b[13]), .CK(clk), .Q(b_whole[13]) );
  DFF_X1 b_reg_reg_12_ ( .D(b[12]), .CK(clk), .Q(b_whole[12]) );
  DFF_X1 b_reg_reg_11_ ( .D(b[11]), .CK(clk), .Q(b_whole[11]) );
  DFF_X1 b_reg_reg_10_ ( .D(b[10]), .CK(clk), .Q(b_whole[10]) );
  DFF_X1 b_reg_reg_9_ ( .D(b[9]), .CK(clk), .Q(b_whole[9]) );
  DFF_X1 b_reg_reg_8_ ( .D(b[8]), .CK(clk), .Q(b_whole[8]) );
  DFF_X1 b_reg_reg_7_ ( .D(b[7]), .CK(clk), .Q(b_whole[7]) );
  DFF_X1 b_reg_reg_6_ ( .D(b[6]), .CK(clk), .Q(b_whole[6]) );
  DFF_X1 b_reg_reg_5_ ( .D(b[5]), .CK(clk), .Q(b_whole[5]) );
  DFF_X1 b_reg_reg_4_ ( .D(b[4]), .CK(clk), .Q(b_whole[4]) );
  DFF_X1 b_reg_reg_3_ ( .D(b[3]), .CK(clk), .Q(b_whole[3]) );
  DFF_X1 b_reg_reg_2_ ( .D(b[2]), .CK(clk), .Q(b_whole[2]) );
  DFF_X1 b_reg_reg_1_ ( .D(b[1]), .CK(clk), .Q(b_whole[1]) );
  DFF_X1 b_reg_reg_0_ ( .D(b[0]), .CK(clk), .Q(b_whole[0]) );
  DFF_X1 result_reg_31_ ( .D(finalSign), .CK(clk), .Q(result[31]) );
  DFF_X1 result_reg_30_ ( .D(outputExponent[7]), .CK(clk), .Q(result[30]) );
  DFF_X1 result_reg_28_ ( .D(outputExponent[5]), .CK(clk), .Q(result[28]) );
  DFF_X1 result_reg_27_ ( .D(outputExponent[4]), .CK(clk), .Q(result[27]) );
  DFF_X1 result_reg_26_ ( .D(outputExponent[3]), .CK(clk), .Q(result[26]) );
  DFF_X1 result_reg_24_ ( .D(outputExponent[1]), .CK(clk), .Q(result[24]) );
  DFF_X1 result_reg_23_ ( .D(outputExponent[0]), .CK(clk), .Q(result[23]) );
  DFF_X1 result_reg_22_ ( .D(normResult[22]), .CK(clk), .Q(result[22]) );
  DFF_X1 result_reg_21_ ( .D(normResult[21]), .CK(clk), .Q(result[21]) );
  DFF_X1 result_reg_20_ ( .D(normResult[20]), .CK(clk), .Q(result[20]) );
  DFF_X1 result_reg_19_ ( .D(normResult[19]), .CK(clk), .Q(result[19]) );
  DFF_X1 result_reg_18_ ( .D(normResult[18]), .CK(clk), .Q(result[18]) );
  DFF_X1 result_reg_17_ ( .D(normResult[17]), .CK(clk), .Q(result[17]) );
  DFF_X1 result_reg_16_ ( .D(normResult[16]), .CK(clk), .Q(result[16]) );
  DFF_X1 result_reg_15_ ( .D(normResult[15]), .CK(clk), .Q(result[15]) );
  DFF_X1 result_reg_14_ ( .D(normResult[14]), .CK(clk), .Q(result[14]) );
  DFF_X1 result_reg_13_ ( .D(normResult[13]), .CK(clk), .Q(result[13]) );
  DFF_X1 result_reg_11_ ( .D(normResult[11]), .CK(clk), .Q(result[11]) );
  DFF_X1 result_reg_9_ ( .D(normResult[9]), .CK(clk), .Q(result[9]) );
  DFF_X1 result_reg_8_ ( .D(normResult[8]), .CK(clk), .Q(result[8]) );
  DFF_X1 result_reg_7_ ( .D(normResult[7]), .CK(clk), .Q(result[7]) );
  DFF_X1 result_reg_6_ ( .D(normResult[6]), .CK(clk), .Q(result[6]) );
  DFF_X1 result_reg_5_ ( .D(normResult[5]), .CK(clk), .Q(result[5]) );
  DFF_X1 result_reg_4_ ( .D(normResult[4]), .CK(clk), .Q(result[4]) );
  DFF_X1 result_reg_3_ ( .D(normResult[3]), .CK(clk), .Q(result[3]) );
  DFF_X1 result_reg_2_ ( .D(normResult[2]), .CK(clk), .Q(result[2]) );
  DFF_X1 result_reg_1_ ( .D(normResult[1]), .CK(clk), .Q(result[1]) );
  DFF_X1 result_reg_0_ ( .D(normResult[0]), .CK(clk), .Q(result[0]) );
  comparator8bit comparator ( .a(a_reg[30:23]), .b(b_reg[30:23]), .f_bigger(
        f_bigger), .diff({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, shiftAmount}) );
  shiftRegister shift ( .a({1'b1, a_whole}), .b({1'b1, b_whole}), .f_bigger(
        n75), .shiftAmount(shiftAmount), .shiftedResult(shiftedResult) );
  Adder24Bit Adder ( .a({1'b1, n97, n98, n99, n101, n102, n103, n104, n105, 
        n106, n107, n108, n109, n110, n89, n90, n91, n92, n93, n94, n95, n96, 
        n100, n111}), .b(shiftedResult), .signFO(signFO), .signSO(signSO), 
        .result(tempResult), .finalSign(finalSign), .cout(cout) );
  Normalize Norm ( .e({n81, n82, n83, n84, n85, n86, n87, n88}), .a(tempResult), .cout(cout), .normExponent(outputExponent), .normResult({
        SYNOPSYS_UNCONNECTED_4, normResult}) );
  DFF_X1 result_reg_12_ ( .D(normResult[12]), .CK(clk), .Q(result[12]) );
  DFF_X1 underflow_reg ( .D(n70), .CK(clk), .Q(underflow) );
  DFF_X1 overflow_reg ( .D(N30), .CK(clk), .Q(overflow) );
  DFF_X1 result_reg_29_ ( .D(outputExponent[6]), .CK(clk), .Q(result[29]) );
  DFF_X1 result_reg_10_ ( .D(normResult[10]), .CK(clk), .Q(result[10]) );
  DFF_X1 result_reg_25_ ( .D(outputExponent[2]), .CK(clk), .Q(result[25]) );
  CLKBUF_X1 U76 ( .A(f_bigger), .Z(n71) );
  BUF_X4 U77 ( .A(n71), .Z(n77) );
  AND4_X1 U78 ( .A1(n76), .A2(n78), .A3(n72), .A4(n73), .ZN(n70) );
  NOR2_X1 U79 ( .A1(outputExponent[2]), .A2(outputExponent[3]), .ZN(n72) );
  NOR2_X1 U80 ( .A1(outputExponent[0]), .A2(outputExponent[1]), .ZN(n73) );
  CLKBUF_X1 U81 ( .A(n75), .Z(n74) );
  BUF_X4 U82 ( .A(f_bigger), .Z(n75) );
  NOR2_X1 U83 ( .A1(outputExponent[6]), .A2(outputExponent[7]), .ZN(n76) );
  NOR2_X1 U84 ( .A1(outputExponent[4]), .A2(outputExponent[5]), .ZN(n78) );
  MUX2_X1 U85 ( .A(b_reg[23]), .B(a_reg[23]), .S(n77), .Z(n88) );
  MUX2_X1 U86 ( .A(b_reg[24]), .B(a_reg[24]), .S(n77), .Z(n87) );
  MUX2_X1 U87 ( .A(b_reg[25]), .B(a_reg[25]), .S(n77), .Z(n86) );
  MUX2_X1 U88 ( .A(b_reg[26]), .B(a_reg[26]), .S(n77), .Z(n85) );
  MUX2_X1 U89 ( .A(b_reg[27]), .B(a_reg[27]), .S(n77), .Z(n84) );
  MUX2_X1 U90 ( .A(b_reg[28]), .B(a_reg[28]), .S(n77), .Z(n83) );
  MUX2_X1 U91 ( .A(b_reg[29]), .B(a_reg[29]), .S(n77), .Z(n82) );
  MUX2_X1 U92 ( .A(b_reg[30]), .B(a_reg[30]), .S(n77), .Z(n81) );
  MUX2_X1 U93 ( .A(a_reg[31]), .B(b_reg[31]), .S(n77), .Z(signSO) );
  MUX2_X1 U94 ( .A(b_reg[31]), .B(a_reg[31]), .S(n74), .Z(signFO) );
  MUX2_X1 U95 ( .A(b_whole[0]), .B(a_whole[0]), .S(n77), .Z(n111) );
  MUX2_X1 U96 ( .A(b_whole[1]), .B(a_whole[1]), .S(n77), .Z(n100) );
  MUX2_X1 U97 ( .A(b_whole[2]), .B(a_whole[2]), .S(n77), .Z(n96) );
  MUX2_X1 U98 ( .A(b_whole[3]), .B(a_whole[3]), .S(n77), .Z(n95) );
  MUX2_X1 U99 ( .A(b_whole[4]), .B(a_whole[4]), .S(n77), .Z(n94) );
  MUX2_X1 U100 ( .A(b_whole[5]), .B(a_whole[5]), .S(n77), .Z(n93) );
  MUX2_X1 U101 ( .A(b_whole[6]), .B(a_whole[6]), .S(n77), .Z(n92) );
  MUX2_X1 U102 ( .A(b_whole[7]), .B(a_whole[7]), .S(n77), .Z(n91) );
  MUX2_X1 U103 ( .A(b_whole[8]), .B(a_whole[8]), .S(n77), .Z(n90) );
  MUX2_X1 U104 ( .A(b_whole[9]), .B(a_whole[9]), .S(n77), .Z(n89) );
  MUX2_X1 U105 ( .A(b_whole[10]), .B(a_whole[10]), .S(n77), .Z(n110) );
  MUX2_X1 U106 ( .A(b_whole[11]), .B(a_whole[11]), .S(n77), .Z(n109) );
  MUX2_X1 U107 ( .A(b_whole[12]), .B(a_whole[12]), .S(n77), .Z(n108) );
  MUX2_X1 U108 ( .A(b_whole[13]), .B(a_whole[13]), .S(n77), .Z(n107) );
  MUX2_X1 U109 ( .A(b_whole[14]), .B(a_whole[14]), .S(n77), .Z(n106) );
  MUX2_X1 U110 ( .A(b_whole[15]), .B(a_whole[15]), .S(n77), .Z(n105) );
  MUX2_X1 U111 ( .A(b_whole[16]), .B(a_whole[16]), .S(n77), .Z(n104) );
  MUX2_X1 U112 ( .A(b_whole[17]), .B(a_whole[17]), .S(n77), .Z(n103) );
  MUX2_X1 U113 ( .A(b_whole[18]), .B(a_whole[18]), .S(n77), .Z(n102) );
  MUX2_X1 U114 ( .A(b_whole[19]), .B(a_whole[19]), .S(n77), .Z(n101) );
  MUX2_X1 U115 ( .A(b_whole[20]), .B(a_whole[20]), .S(n77), .Z(n99) );
  MUX2_X1 U116 ( .A(b_whole[21]), .B(a_whole[21]), .S(n77), .Z(n98) );
  MUX2_X1 U117 ( .A(b_whole[22]), .B(a_whole[22]), .S(n77), .Z(n97) );
  NAND4_X1 U118 ( .A1(outputExponent[3]), .A2(outputExponent[2]), .A3(
        outputExponent[1]), .A4(outputExponent[0]), .ZN(n80) );
  NAND4_X1 U119 ( .A1(outputExponent[6]), .A2(outputExponent[4]), .A3(
        outputExponent[5]), .A4(outputExponent[7]), .ZN(n79) );
  NOR2_X1 U120 ( .A1(n79), .A2(n80), .ZN(N30) );
endmodule

