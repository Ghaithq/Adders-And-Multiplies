
module FPMultiplier_DW01_add_1 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [7:2] carry;

  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module FPMultiplier_DW_mult_uns_0 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n174, n175, n177, n178, n180, n181, n182, n183, n184,
         n185, n186, n187, n189, n190, n191, n192, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n207, n208, n209,
         n210, n211, n212, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n231, n232, n233,
         n234, n235, n236, n237, n238, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n555, n556, n557, n558, n559, n560, n561, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n665, n667, n669,
         n671, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n875, n876,
         n877, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337;

  FA_X1 U128 ( .A(n178), .B(n180), .CI(n128), .CO(n127), .S(product[45]) );
  FA_X1 U130 ( .A(n185), .B(n189), .CI(n130), .CO(n129), .S(product[43]) );
  FA_X1 U132 ( .A(n195), .B(n200), .CI(n132), .CO(n131), .S(product[41]) );
  FA_X1 U134 ( .A(n208), .B(n214), .CI(n134), .CO(n133), .S(product[39]) );
  FA_X1 U136 ( .A(n223), .B(n231), .CI(n136), .CO(n135), .S(product[37]) );
  FA_X1 U139 ( .A(n251), .B(n261), .CI(n139), .CO(n138), .S(product[34]) );
  FA_X1 U143 ( .A(n298), .B(n310), .CI(n143), .CO(n142), .S(product[30]) );
  FA_X1 U147 ( .A(n353), .B(n366), .CI(n147), .CO(n146), .S(product[26]) );
  FA_X1 U150 ( .A(n877), .B(n395), .CI(n150), .CO(n149), .S(product[23]) );
  FA_X1 U175 ( .A(n1839), .B(b[22]), .CI(n687), .CO(n174), .S(n175) );
  FA_X1 U177 ( .A(n182), .B(n1839), .CI(n688), .CO(n177), .S(n178) );
  FA_X1 U179 ( .A(n689), .B(n183), .CI(n186), .CO(n180), .S(n181) );
  FA_X1 U180 ( .A(b[19]), .B(n1762), .CI(b[20]), .CO(n182), .S(n183) );
  FA_X1 U181 ( .A(n713), .B(n690), .CI(n187), .CO(n184), .S(n185) );
  FA_X1 U182 ( .A(n1842), .B(b[18]), .CI(n191), .CO(n186), .S(n187) );
  FA_X1 U184 ( .A(n192), .B(n196), .CI(n714), .CO(n189), .S(n190) );
  FA_X1 U185 ( .A(n198), .B(n1844), .CI(n691), .CO(n191), .S(n192) );
  FA_X1 U187 ( .A(n715), .B(n197), .CI(n202), .CO(n194), .S(n195) );
  FA_X1 U188 ( .A(n204), .B(n199), .CI(n692), .CO(n196), .S(n197) );
  FA_X1 U189 ( .A(b[17]), .B(n1764), .CI(b[15]), .CO(n198), .S(n199) );
  FA_X1 U190 ( .A(n740), .B(n716), .CI(n203), .CO(n200), .S(n201) );
  FA_X1 U191 ( .A(n205), .B(n211), .CI(n209), .CO(n202), .S(n203) );
  FA_X1 U192 ( .A(n1848), .B(b[16]), .CI(n693), .CO(n204), .S(n205) );
  FA_X1 U194 ( .A(n210), .B(n216), .CI(n741), .CO(n207), .S(n208) );
  FA_X1 U195 ( .A(n212), .B(n218), .CI(n717), .CO(n209), .S(n210) );
  FA_X1 U196 ( .A(n220), .B(n1848), .CI(n694), .CO(n211), .S(n212) );
  FA_X1 U198 ( .A(n742), .B(n217), .CI(n224), .CO(n214), .S(n215) );
  FA_X1 U199 ( .A(n226), .B(n219), .CI(n718), .CO(n216), .S(n217) );
  FA_X1 U200 ( .A(n228), .B(n221), .CI(n695), .CO(n218), .S(n219) );
  FA_X1 U201 ( .A(b[13]), .B(n1766), .CI(b[14]), .CO(n220), .S(n221) );
  FA_X1 U202 ( .A(n767), .B(n743), .CI(n225), .CO(n222), .S(n223) );
  FA_X1 U203 ( .A(n227), .B(n235), .CI(n233), .CO(n224), .S(n225) );
  FA_X1 U204 ( .A(n229), .B(n696), .CI(n719), .CO(n226), .S(n227) );
  FA_X1 U205 ( .A(n1852), .B(b[12]), .CI(n237), .CO(n228), .S(n229) );
  FA_X1 U207 ( .A(n234), .B(n242), .CI(n768), .CO(n231), .S(n232) );
  FA_X1 U208 ( .A(n236), .B(n244), .CI(n744), .CO(n233), .S(n234) );
  FA_X1 U209 ( .A(n238), .B(n246), .CI(n720), .CO(n235), .S(n236) );
  FA_X1 U210 ( .A(n248), .B(n1854), .CI(n697), .CO(n237), .S(n238) );
  FA_X1 U212 ( .A(n769), .B(n243), .CI(n252), .CO(n240), .S(n241) );
  FA_X1 U213 ( .A(n254), .B(n245), .CI(n745), .CO(n242), .S(n243) );
  FA_X1 U214 ( .A(n721), .B(n247), .CI(n256), .CO(n244), .S(n245) );
  FA_X1 U215 ( .A(n258), .B(n249), .CI(n698), .CO(n246), .S(n247) );
  FA_X1 U216 ( .A(b[11]), .B(n1768), .CI(b[9]), .CO(n248), .S(n249) );
  FA_X1 U217 ( .A(n794), .B(n770), .CI(n253), .CO(n250), .S(n251) );
  FA_X1 U218 ( .A(n255), .B(n265), .CI(n263), .CO(n252), .S(n253) );
  FA_X1 U219 ( .A(n257), .B(n722), .CI(n746), .CO(n254), .S(n255) );
  FA_X1 U220 ( .A(n259), .B(n269), .CI(n267), .CO(n256), .S(n257) );
  FA_X1 U221 ( .A(n1860), .B(b[10]), .CI(n699), .CO(n258), .S(n259) );
  FA_X1 U223 ( .A(n264), .B(n274), .CI(n795), .CO(n261), .S(n262) );
  FA_X1 U224 ( .A(n266), .B(n276), .CI(n771), .CO(n263), .S(n264) );
  FA_X1 U225 ( .A(n268), .B(n278), .CI(n747), .CO(n265), .S(n266) );
  FA_X1 U226 ( .A(n270), .B(n280), .CI(n723), .CO(n267), .S(n268) );
  FA_X1 U227 ( .A(n282), .B(n1860), .CI(n700), .CO(n269), .S(n270) );
  FA_X1 U229 ( .A(n796), .B(n275), .CI(n286), .CO(n272), .S(n273) );
  FA_X1 U230 ( .A(n288), .B(n277), .CI(n772), .CO(n274), .S(n275) );
  FA_X1 U231 ( .A(n748), .B(n279), .CI(n290), .CO(n276), .S(n277) );
  FA_X1 U232 ( .A(n292), .B(n281), .CI(n724), .CO(n278), .S(n279) );
  FA_X1 U233 ( .A(n701), .B(n283), .CI(n294), .CO(n280), .S(n281) );
  FA_X1 U234 ( .A(b[7]), .B(n1770), .CI(b[8]), .CO(n282), .S(n283) );
  FA_X1 U235 ( .A(n821), .B(n797), .CI(n287), .CO(n284), .S(n285) );
  FA_X1 U236 ( .A(n289), .B(n301), .CI(n299), .CO(n286), .S(n287) );
  FA_X1 U237 ( .A(n291), .B(n749), .CI(n773), .CO(n288), .S(n289) );
  FA_X1 U238 ( .A(n293), .B(n725), .CI(n303), .CO(n290), .S(n291) );
  FA_X1 U239 ( .A(n295), .B(n702), .CI(n305), .CO(n292), .S(n293) );
  FA_X1 U240 ( .A(n1864), .B(b[6]), .CI(n307), .CO(n294), .S(n295) );
  FA_X1 U242 ( .A(n300), .B(n312), .CI(n822), .CO(n297), .S(n298) );
  FA_X1 U243 ( .A(n302), .B(n314), .CI(n798), .CO(n299), .S(n300) );
  FA_X1 U244 ( .A(n304), .B(n316), .CI(n774), .CO(n301), .S(n302) );
  FA_X1 U245 ( .A(n306), .B(n318), .CI(n750), .CO(n303), .S(n304) );
  FA_X1 U246 ( .A(n308), .B(n320), .CI(n726), .CO(n305), .S(n306) );
  FA_X1 U247 ( .A(n322), .B(n1866), .CI(n703), .CO(n307), .S(n308) );
  FA_X1 U249 ( .A(n823), .B(n313), .CI(n326), .CO(n310), .S(n311) );
  FA_X1 U250 ( .A(n328), .B(n315), .CI(n799), .CO(n312), .S(n313) );
  FA_X1 U251 ( .A(n330), .B(n317), .CI(n775), .CO(n314), .S(n315) );
  FA_X1 U252 ( .A(n332), .B(n319), .CI(n751), .CO(n316), .S(n317) );
  FA_X1 U253 ( .A(n334), .B(n321), .CI(n727), .CO(n318), .S(n319) );
  FA_X1 U254 ( .A(n336), .B(n323), .CI(n704), .CO(n320), .S(n321) );
  FA_X1 U255 ( .A(n1496), .B(n1772), .CI(b[5]), .CO(n322), .S(n323) );
  FA_X1 U256 ( .A(n848), .B(n824), .CI(n327), .CO(n324), .S(n325) );
  FA_X1 U257 ( .A(n329), .B(n342), .CI(n340), .CO(n326), .S(n327) );
  FA_X1 U258 ( .A(n331), .B(n776), .CI(n800), .CO(n328), .S(n329) );
  FA_X1 U259 ( .A(n333), .B(n752), .CI(n344), .CO(n330), .S(n331) );
  FA_X1 U260 ( .A(n335), .B(n728), .CI(n346), .CO(n332), .S(n333) );
  FA_X1 U261 ( .A(n337), .B(n705), .CI(n348), .CO(n334), .S(n335) );
  FA_X1 U262 ( .A(b[4]), .B(n1482), .CI(n350), .CO(n336), .S(n337) );
  FA_X1 U263 ( .A(n341), .B(n825), .CI(n849), .CO(n338), .S(n339) );
  FA_X1 U264 ( .A(n343), .B(n356), .CI(n354), .CO(n340), .S(n341) );
  FA_X1 U265 ( .A(n345), .B(n777), .CI(n801), .CO(n342), .S(n343) );
  FA_X1 U266 ( .A(n347), .B(n360), .CI(n358), .CO(n344), .S(n345) );
  FA_X1 U267 ( .A(n349), .B(n729), .CI(n753), .CO(n346), .S(n347) );
  FA_X1 U268 ( .A(n351), .B(n364), .CI(n362), .CO(n348), .S(n349) );
  FA_X1 U269 ( .A(b[3]), .B(n1482), .CI(n706), .CO(n350), .S(n351) );
  FA_X1 U270 ( .A(n355), .B(n368), .CI(n850), .CO(n352), .S(n353) );
  FA_X1 U271 ( .A(n357), .B(n370), .CI(n826), .CO(n354), .S(n355) );
  FA_X1 U272 ( .A(n359), .B(n372), .CI(n802), .CO(n356), .S(n357) );
  FA_X1 U273 ( .A(n361), .B(n374), .CI(n778), .CO(n358), .S(n359) );
  FA_X1 U274 ( .A(n363), .B(n376), .CI(n754), .CO(n360), .S(n361) );
  FA_X1 U275 ( .A(n365), .B(n378), .CI(n730), .CO(n362), .S(n363) );
  FA_X1 U276 ( .A(n1649), .B(n1482), .CI(n707), .CO(n364), .S(n365) );
  FA_X1 U277 ( .A(n851), .B(n369), .CI(n875), .CO(n366), .S(n367) );
  FA_X1 U278 ( .A(n827), .B(n371), .CI(n382), .CO(n368), .S(n369) );
  FA_X1 U279 ( .A(n803), .B(n373), .CI(n384), .CO(n370), .S(n371) );
  FA_X1 U280 ( .A(n779), .B(n375), .CI(n386), .CO(n372), .S(n373) );
  FA_X1 U281 ( .A(n755), .B(n377), .CI(n388), .CO(n374), .S(n375) );
  FA_X1 U282 ( .A(n731), .B(n379), .CI(n390), .CO(n376), .S(n377) );
  FA_X1 U283 ( .A(n708), .B(n1745), .CI(n392), .CO(n378), .S(n379) );
  FA_X1 U284 ( .A(n852), .B(n383), .CI(n394), .CO(n380), .S(n381) );
  FA_X1 U285 ( .A(n828), .B(n385), .CI(n396), .CO(n382), .S(n383) );
  FA_X1 U286 ( .A(n804), .B(n387), .CI(n398), .CO(n384), .S(n385) );
  FA_X1 U287 ( .A(n780), .B(n389), .CI(n400), .CO(n386), .S(n387) );
  FA_X1 U288 ( .A(n756), .B(n391), .CI(n402), .CO(n388), .S(n389) );
  FA_X1 U289 ( .A(n732), .B(n393), .CI(n404), .CO(n390), .S(n391) );
  FA_X1 U290 ( .A(n406), .B(n1716), .CI(n709), .CO(n392), .S(n393) );
  FA_X1 U293 ( .A(n805), .B(n401), .CI(n412), .CO(n398), .S(n399) );
  FA_X1 U294 ( .A(n781), .B(n403), .CI(n414), .CO(n400), .S(n401) );
  FA_X1 U295 ( .A(n757), .B(n405), .CI(n416), .CO(n402), .S(n403) );
  FA_X1 U296 ( .A(n733), .B(n407), .CI(n418), .CO(n404), .S(n405) );
  HA_X1 U297 ( .A(n420), .B(n710), .CO(n406), .S(n407) );
  FA_X1 U298 ( .A(n854), .B(n411), .CI(n422), .CO(n408), .S(n409) );
  FA_X1 U300 ( .A(n806), .B(n415), .CI(n426), .CO(n412), .S(n413) );
  FA_X1 U301 ( .A(n782), .B(n417), .CI(n428), .CO(n414), .S(n415) );
  FA_X1 U302 ( .A(n758), .B(n419), .CI(n430), .CO(n416), .S(n417) );
  FA_X1 U303 ( .A(n734), .B(n421), .CI(n432), .CO(n418), .S(n419) );
  HA_X1 U304 ( .A(n711), .B(n434), .CO(n420), .S(n421) );
  FA_X1 U306 ( .A(n831), .B(n427), .CI(n438), .CO(n424), .S(n425) );
  FA_X1 U307 ( .A(n807), .B(n429), .CI(n440), .CO(n426), .S(n427) );
  FA_X1 U308 ( .A(n783), .B(n431), .CI(n442), .CO(n428), .S(n429) );
  FA_X1 U309 ( .A(n759), .B(n433), .CI(n444), .CO(n430), .S(n431) );
  FA_X1 U310 ( .A(n735), .B(n1798), .CI(n446), .CO(n432), .S(n433) );
  FA_X1 U312 ( .A(n856), .B(n439), .CI(n448), .CO(n436), .S(n437) );
  FA_X1 U314 ( .A(n808), .B(n443), .CI(n452), .CO(n440), .S(n441) );
  FA_X1 U315 ( .A(n784), .B(n445), .CI(n454), .CO(n442), .S(n443) );
  FA_X1 U316 ( .A(n760), .B(n447), .CI(n456), .CO(n444), .S(n445) );
  HA_X1 U317 ( .A(n458), .B(n736), .CO(n446), .S(n447) );
  FA_X1 U319 ( .A(n833), .B(n453), .CI(n462), .CO(n450), .S(n451) );
  FA_X1 U320 ( .A(n809), .B(n455), .CI(n464), .CO(n452), .S(n453) );
  FA_X1 U321 ( .A(n785), .B(n457), .CI(n466), .CO(n454), .S(n455) );
  FA_X1 U322 ( .A(n761), .B(n459), .CI(n468), .CO(n456), .S(n457) );
  HA_X1 U323 ( .A(n470), .B(n737), .CO(n458), .S(n459) );
  FA_X1 U325 ( .A(n834), .B(n465), .CI(n474), .CO(n462), .S(n463) );
  FA_X1 U326 ( .A(n810), .B(n467), .CI(n476), .CO(n464), .S(n465) );
  FA_X1 U327 ( .A(n786), .B(n469), .CI(n478), .CO(n466), .S(n467) );
  FA_X1 U328 ( .A(n762), .B(n471), .CI(n480), .CO(n468), .S(n469) );
  HA_X1 U329 ( .A(n738), .B(a[20]), .CO(n470), .S(n471) );
  FA_X1 U331 ( .A(n835), .B(n477), .CI(n484), .CO(n474), .S(n475) );
  FA_X1 U332 ( .A(n811), .B(n479), .CI(n486), .CO(n476), .S(n477) );
  FA_X1 U333 ( .A(n787), .B(n481), .CI(n488), .CO(n478), .S(n479) );
  HA_X1 U334 ( .A(n490), .B(n763), .CO(n480), .S(n481) );
  FA_X1 U336 ( .A(n836), .B(n487), .CI(n494), .CO(n484), .S(n485) );
  FA_X1 U337 ( .A(n812), .B(n489), .CI(n496), .CO(n486), .S(n487) );
  FA_X1 U338 ( .A(n788), .B(n491), .CI(n498), .CO(n488), .S(n489) );
  HA_X1 U339 ( .A(n500), .B(n764), .CO(n490), .S(n491) );
  FA_X1 U340 ( .A(n861), .B(n495), .CI(n502), .CO(n492), .S(n493) );
  FA_X1 U341 ( .A(n837), .B(n497), .CI(n504), .CO(n494), .S(n495) );
  FA_X1 U342 ( .A(n813), .B(n499), .CI(n506), .CO(n496), .S(n497) );
  FA_X1 U343 ( .A(n789), .B(n501), .CI(n508), .CO(n498), .S(n499) );
  HA_X1 U344 ( .A(n765), .B(a[17]), .CO(n500), .S(n501) );
  FA_X1 U347 ( .A(n814), .B(n509), .CI(n514), .CO(n506), .S(n507) );
  HA_X1 U348 ( .A(n516), .B(n790), .CO(n508), .S(n509) );
  FA_X1 U350 ( .A(n839), .B(n515), .CI(n520), .CO(n512), .S(n513) );
  FA_X1 U351 ( .A(n815), .B(n517), .CI(n522), .CO(n514), .S(n515) );
  HA_X1 U352 ( .A(n524), .B(n791), .CO(n516), .S(n517) );
  FA_X1 U354 ( .A(n840), .B(n523), .CI(n528), .CO(n520), .S(n521) );
  FA_X1 U355 ( .A(n816), .B(n525), .CI(n530), .CO(n522), .S(n523) );
  HA_X1 U356 ( .A(n792), .B(a[14]), .CO(n524), .S(n525) );
  FA_X1 U358 ( .A(n841), .B(n531), .CI(n534), .CO(n528), .S(n529) );
  HA_X1 U359 ( .A(n536), .B(n817), .CO(n530), .S(n531) );
  FA_X1 U360 ( .A(n866), .B(n535), .CI(n538), .CO(n532), .S(n533) );
  FA_X1 U361 ( .A(n842), .B(n537), .CI(n540), .CO(n534), .S(n535) );
  HA_X1 U362 ( .A(n542), .B(n818), .CO(n536), .S(n537) );
  HA_X1 U365 ( .A(n819), .B(a[11]), .CO(n542), .S(n543) );
  FA_X1 U366 ( .A(n868), .B(n547), .CI(n548), .CO(n544), .S(n545) );
  HA_X1 U367 ( .A(n550), .B(n844), .CO(n546), .S(n547) );
  FA_X1 U368 ( .A(n869), .B(n551), .CI(n552), .CO(n548), .S(n549) );
  HA_X1 U369 ( .A(n1478), .B(n845), .CO(n550), .S(n551) );
  FA_X1 U370 ( .A(n870), .B(n556), .CI(n555), .CO(n552), .S(n553) );
  HA_X1 U372 ( .A(n558), .B(n871), .CO(n556), .S(n557) );
  HA_X1 U373 ( .A(n560), .B(n872), .CO(n558), .S(n559) );
  HA_X1 U374 ( .A(n873), .B(a[5]), .CO(n560), .S(n561) );
  FA_X1 U1163 ( .A(b[21]), .B(b[22]), .CI(n642), .CO(n641), .S(n665) );
  FA_X1 U1165 ( .A(b[19]), .B(b[20]), .CI(n644), .CO(n643), .S(n667) );
  FA_X1 U1167 ( .A(b[17]), .B(b[18]), .CI(n646), .CO(n645), .S(n669) );
  FA_X1 U1169 ( .A(b[15]), .B(b[16]), .CI(n648), .CO(n647), .S(n671) );
  FA_X1 U1171 ( .A(b[13]), .B(b[14]), .CI(n650), .CO(n649), .S(n673) );
  FA_X1 U1173 ( .A(b[11]), .B(b[12]), .CI(n652), .CO(n651), .S(n675) );
  FA_X1 U1175 ( .A(b[9]), .B(b[10]), .CI(n654), .CO(n653), .S(n677) );
  FA_X1 U1177 ( .A(b[7]), .B(b[8]), .CI(n656), .CO(n655), .S(n679) );
  FA_X1 U1179 ( .A(b[5]), .B(b[6]), .CI(n658), .CO(n657), .S(n681) );
  FA_X1 U1180 ( .A(b[4]), .B(b[5]), .CI(n659), .CO(n658), .S(n682) );
  FA_X1 U1182 ( .A(b[2]), .B(b[3]), .CI(n661), .CO(n660), .S(n684) );
  INV_X2 U1188 ( .A(n1883), .ZN(n1829) );
  INV_X2 U1189 ( .A(n1484), .ZN(n1895) );
  BUF_X2 U1190 ( .A(n1944), .Z(n1783) );
  AND3_X1 U1191 ( .A1(n1524), .A2(n1525), .A3(n1526), .ZN(n2327) );
  AND3_X1 U1192 ( .A1(n1679), .A2(n1680), .A3(n1681), .ZN(n2311) );
  OAI221_X1 U1193 ( .B1(n1848), .B2(n1483), .C1(n1777), .C2(n1634), .A(n1925), 
        .ZN(n1924) );
  AOI221_X1 U1194 ( .B1(n2171), .B2(b[22]), .C1(n1620), .C2(n1497), .A(n2212), 
        .ZN(n2211) );
  OAI221_X1 U1195 ( .B1(n1844), .B2(n1947), .C1(n1840), .C2(n1783), .A(n1985), 
        .ZN(n1984) );
  NAND2_X1 U1196 ( .A1(n2335), .A2(a[0]), .ZN(n1883) );
  BUF_X2 U1197 ( .A(n1890), .Z(n1777) );
  AOI221_X1 U1198 ( .B1(n1793), .B2(b[22]), .C1(n2223), .C2(n1497), .A(n2245), 
        .ZN(n690) );
  INV_X1 U1199 ( .A(n1622), .ZN(n1471) );
  INV_X1 U1200 ( .A(n1622), .ZN(n1785) );
  OR2_X2 U1201 ( .A1(n1479), .A2(n1996), .ZN(n1622) );
  AND2_X1 U1202 ( .A1(n1816), .A2(n2104), .ZN(n1472) );
  OR2_X1 U1203 ( .A1(n1625), .A2(n1941), .ZN(n1473) );
  XOR2_X1 U1204 ( .A(n1573), .B(n1618), .Z(n1474) );
  XNOR2_X1 U1205 ( .A(n1512), .B(n1507), .ZN(n1475) );
  XOR2_X1 U1206 ( .A(n1571), .B(n1617), .Z(n1476) );
  XNOR2_X1 U1207 ( .A(n492), .B(n1593), .ZN(n1477) );
  AND2_X1 U1208 ( .A1(n846), .A2(a[8]), .ZN(n1478) );
  XNOR2_X1 U1209 ( .A(a[6]), .B(n1773), .ZN(n1479) );
  NAND2_X1 U1210 ( .A1(n1635), .A2(n1636), .ZN(n1480) );
  OR2_X1 U1211 ( .A1(n1700), .A2(n1701), .ZN(n1481) );
  NOR2_X2 U1212 ( .A1(n1834), .A2(n2335), .ZN(n2294) );
  XNOR2_X1 U1213 ( .A(a[9]), .B(a[8]), .ZN(n2049) );
  AND3_X1 U1214 ( .A1(n1676), .A2(n1677), .A3(n1678), .ZN(n2278) );
  CLKBUF_X1 U1215 ( .A(a[2]), .Z(n1482) );
  INV_X1 U1216 ( .A(n1827), .ZN(n1483) );
  NAND3_X1 U1217 ( .A1(n1647), .A2(n1732), .A3(n1941), .ZN(n1893) );
  OAI221_X1 U1218 ( .B1(n1852), .B2(n1483), .C1(n1777), .C2(n1632), .A(n1921), 
        .ZN(n1920) );
  XOR2_X2 U1219 ( .A(n1587), .B(n1633), .Z(n1632) );
  XNOR2_X2 U1220 ( .A(n1506), .B(n1667), .ZN(n1634) );
  NAND2_X1 U1221 ( .A1(n1624), .A2(n1625), .ZN(n1484) );
  INV_X1 U1222 ( .A(n667), .ZN(n1485) );
  INV_X1 U1223 ( .A(n667), .ZN(n1840) );
  CLKBUF_X1 U1224 ( .A(n1630), .Z(n1486) );
  CLKBUF_X1 U1225 ( .A(n645), .Z(n1487) );
  XOR2_X1 U1226 ( .A(a[6]), .B(n1773), .Z(n1488) );
  CLKBUF_X1 U1227 ( .A(n1491), .Z(n1489) );
  INV_X1 U1228 ( .A(n1588), .ZN(n1490) );
  INV_X1 U1229 ( .A(n1588), .ZN(n1949) );
  NAND3_X1 U1230 ( .A1(n1726), .A2(n1725), .A3(n1727), .ZN(n1491) );
  INV_X1 U1231 ( .A(n2218), .ZN(n1492) );
  CLKBUF_X1 U1232 ( .A(n1486), .Z(n1493) );
  CLKBUF_X1 U1233 ( .A(n1628), .Z(n1494) );
  INV_X1 U1234 ( .A(n669), .ZN(n1495) );
  AND3_X1 U1235 ( .A1(n1580), .A2(n1581), .A3(n1582), .ZN(n2271) );
  CLKBUF_X1 U1236 ( .A(n1831), .Z(n1496) );
  INV_X1 U1237 ( .A(a[2]), .ZN(n1831) );
  INV_X1 U1238 ( .A(n1837), .ZN(n1497) );
  XOR2_X1 U1239 ( .A(n441), .B(n832), .Z(n1498) );
  XOR2_X1 U1240 ( .A(n450), .B(n1498), .Z(n439) );
  NAND2_X1 U1241 ( .A1(n450), .A2(n441), .ZN(n1499) );
  NAND2_X1 U1242 ( .A1(n450), .A2(n832), .ZN(n1500) );
  NAND2_X1 U1243 ( .A1(n441), .A2(n832), .ZN(n1501) );
  NAND3_X1 U1244 ( .A1(n1499), .A2(n1500), .A3(n1501), .ZN(n438) );
  XOR2_X1 U1245 ( .A(n543), .B(n843), .Z(n1502) );
  XOR2_X1 U1246 ( .A(n546), .B(n1502), .Z(n541) );
  NAND2_X1 U1247 ( .A1(n546), .A2(n543), .ZN(n1503) );
  NAND2_X1 U1248 ( .A1(n546), .A2(n843), .ZN(n1504) );
  NAND2_X1 U1249 ( .A1(n543), .A2(n843), .ZN(n1505) );
  NAND3_X1 U1250 ( .A1(n1503), .A2(n1504), .A3(n1505), .ZN(n540) );
  XNOR2_X1 U1251 ( .A(n1912), .B(n1773), .ZN(n862) );
  CLKBUF_X1 U1252 ( .A(n647), .Z(n1506) );
  XOR2_X1 U1253 ( .A(n505), .B(n862), .Z(n1507) );
  NAND2_X1 U1254 ( .A1(n1511), .A2(n505), .ZN(n1508) );
  NAND2_X1 U1255 ( .A1(n510), .A2(n862), .ZN(n1509) );
  NAND2_X1 U1256 ( .A1(n505), .A2(n862), .ZN(n1510) );
  NAND3_X1 U1257 ( .A1(n1508), .A2(n1509), .A3(n1510), .ZN(n502) );
  NAND3_X1 U1258 ( .A1(n1641), .A2(n1642), .A3(n1643), .ZN(n1511) );
  NAND3_X1 U1259 ( .A1(n1641), .A2(n1642), .A3(n1643), .ZN(n1512) );
  AND3_X2 U1260 ( .A1(n1606), .A2(n1607), .A3(n1608), .ZN(n2263) );
  CLKBUF_X1 U1261 ( .A(n660), .Z(n1513) );
  CLKBUF_X1 U1262 ( .A(n651), .Z(n1514) );
  CLKBUF_X1 U1263 ( .A(n653), .Z(n1515) );
  CLKBUF_X1 U1264 ( .A(n146), .Z(n1516) );
  OR2_X2 U1265 ( .A1(n1993), .A2(n1488), .ZN(n1588) );
  CLKBUF_X1 U1266 ( .A(n1944), .Z(n1782) );
  XNOR2_X1 U1267 ( .A(n1517), .B(n410), .ZN(n397) );
  XNOR2_X1 U1268 ( .A(n829), .B(n399), .ZN(n1517) );
  XNOR2_X1 U1269 ( .A(n408), .B(n1518), .ZN(n395) );
  XNOR2_X1 U1270 ( .A(n397), .B(n853), .ZN(n1518) );
  CLKBUF_X1 U1271 ( .A(b[1]), .Z(n1519) );
  CLKBUF_X1 U1272 ( .A(n1542), .Z(n1520) );
  CLKBUF_X1 U1273 ( .A(n149), .Z(n1521) );
  CLKBUF_X1 U1274 ( .A(n1543), .Z(n1522) );
  NAND3_X1 U1275 ( .A1(n1536), .A2(n1537), .A3(n1538), .ZN(n1523) );
  NOR2_X1 U1276 ( .A1(n2266), .A2(n1481), .ZN(n2265) );
  CLKBUF_X1 U1277 ( .A(n657), .Z(n1601) );
  NAND2_X1 U1278 ( .A1(n2331), .A2(n2332), .ZN(n1524) );
  NAND2_X1 U1279 ( .A1(n2331), .A2(n561), .ZN(n1525) );
  NAND2_X1 U1280 ( .A1(n561), .A2(n2332), .ZN(n1526) );
  AND3_X2 U1281 ( .A1(n1638), .A2(n1639), .A3(n1640), .ZN(n2286) );
  XOR2_X1 U1282 ( .A(n324), .B(n311), .Z(n1527) );
  XOR2_X1 U1283 ( .A(n1532), .B(n1527), .Z(product[29]) );
  NAND2_X1 U1284 ( .A1(n1531), .A2(n324), .ZN(n1528) );
  NAND2_X1 U1285 ( .A1(n144), .A2(n311), .ZN(n1529) );
  NAND2_X1 U1286 ( .A1(n324), .A2(n311), .ZN(n1530) );
  NAND3_X1 U1287 ( .A1(n1528), .A2(n1529), .A3(n1530), .ZN(n143) );
  NAND3_X1 U1288 ( .A1(n1687), .A2(n1686), .A3(n1688), .ZN(n1531) );
  NAND3_X1 U1289 ( .A1(n1687), .A2(n1686), .A3(n1688), .ZN(n1532) );
  CLKBUF_X1 U1290 ( .A(n655), .Z(n1533) );
  CLKBUF_X1 U1291 ( .A(n1519), .Z(n1534) );
  XOR2_X1 U1292 ( .A(n339), .B(n352), .Z(n1535) );
  XOR2_X1 U1293 ( .A(n1516), .B(n1535), .Z(product[27]) );
  NAND2_X1 U1294 ( .A1(n146), .A2(n339), .ZN(n1536) );
  NAND2_X1 U1295 ( .A1(n146), .A2(n352), .ZN(n1537) );
  NAND2_X1 U1296 ( .A1(n339), .A2(n352), .ZN(n1538) );
  NAND3_X1 U1297 ( .A1(n1537), .A2(n1536), .A3(n1538), .ZN(n145) );
  CLKBUF_X1 U1298 ( .A(n133), .Z(n1539) );
  CLKBUF_X1 U1299 ( .A(n129), .Z(n1540) );
  CLKBUF_X1 U1300 ( .A(n142), .Z(n1541) );
  NAND3_X1 U1301 ( .A1(n1697), .A2(n1698), .A3(n1699), .ZN(n1542) );
  NAND3_X1 U1302 ( .A1(n1709), .A2(n1710), .A3(n1711), .ZN(n1543) );
  AND2_X1 U1303 ( .A1(b[0]), .A2(n1534), .ZN(n1545) );
  AND2_X1 U1304 ( .A1(b[1]), .A2(b[0]), .ZN(n1544) );
  AND2_X1 U1305 ( .A1(b[0]), .A2(b[1]), .ZN(n1648) );
  XOR2_X1 U1306 ( .A(n830), .B(n413), .Z(n1546) );
  XOR2_X1 U1307 ( .A(n1546), .B(n424), .Z(n411) );
  NAND2_X1 U1308 ( .A1(n830), .A2(n413), .ZN(n1547) );
  NAND2_X1 U1309 ( .A1(n830), .A2(n424), .ZN(n1548) );
  NAND2_X1 U1310 ( .A1(n413), .A2(n424), .ZN(n1549) );
  NAND3_X1 U1311 ( .A1(n1547), .A2(n1548), .A3(n1549), .ZN(n410) );
  NAND2_X1 U1312 ( .A1(n829), .A2(n399), .ZN(n1550) );
  NAND2_X1 U1313 ( .A1(n829), .A2(n410), .ZN(n1551) );
  NAND2_X1 U1314 ( .A1(n399), .A2(n410), .ZN(n1552) );
  NAND3_X1 U1315 ( .A1(n1550), .A2(n1551), .A3(n1552), .ZN(n396) );
  XOR2_X1 U1316 ( .A(n507), .B(n838), .Z(n1553) );
  XOR2_X1 U1317 ( .A(n512), .B(n1553), .Z(n505) );
  NAND2_X1 U1318 ( .A1(n512), .A2(n507), .ZN(n1554) );
  NAND2_X1 U1319 ( .A1(n512), .A2(n838), .ZN(n1555) );
  NAND2_X1 U1320 ( .A1(n507), .A2(n838), .ZN(n1556) );
  NAND3_X1 U1321 ( .A1(n1554), .A2(n1555), .A3(n1556), .ZN(n504) );
  XOR2_X1 U1322 ( .A(b[2]), .B(n1519), .Z(n1557) );
  XOR2_X1 U1323 ( .A(n1545), .B(n1557), .Z(n685) );
  NAND2_X1 U1324 ( .A1(n1544), .A2(b[2]), .ZN(n1558) );
  NAND2_X1 U1325 ( .A1(n1648), .A2(b[1]), .ZN(n1559) );
  NAND2_X1 U1326 ( .A1(b[1]), .A2(b[2]), .ZN(n1560) );
  NAND3_X1 U1327 ( .A1(n1558), .A2(n1559), .A3(n1560), .ZN(n661) );
  XOR2_X1 U1328 ( .A(b[13]), .B(b[12]), .Z(n1561) );
  XOR2_X1 U1329 ( .A(n1514), .B(n1561), .Z(n674) );
  NAND2_X1 U1330 ( .A1(n651), .A2(b[13]), .ZN(n1562) );
  NAND2_X1 U1331 ( .A1(n651), .A2(b[12]), .ZN(n1563) );
  NAND2_X1 U1332 ( .A1(b[13]), .A2(b[12]), .ZN(n1564) );
  NAND3_X1 U1333 ( .A1(n1562), .A2(n1563), .A3(n1564), .ZN(n650) );
  NAND2_X1 U1334 ( .A1(n408), .A2(n397), .ZN(n1565) );
  NAND2_X1 U1335 ( .A1(n408), .A2(n853), .ZN(n1566) );
  NAND2_X1 U1336 ( .A1(n397), .A2(n853), .ZN(n1567) );
  NAND3_X1 U1337 ( .A1(n1565), .A2(n1566), .A3(n1567), .ZN(n394) );
  NAND3_X1 U1338 ( .A1(n1594), .A2(n1595), .A3(n1596), .ZN(n1568) );
  NAND3_X1 U1339 ( .A1(n1594), .A2(n1595), .A3(n1596), .ZN(n1569) );
  NAND3_X1 U1340 ( .A1(n1759), .A2(n1760), .A3(n1761), .ZN(n1570) );
  NAND3_X1 U1341 ( .A1(n1759), .A2(n1760), .A3(n1761), .ZN(n1571) );
  NAND3_X1 U1342 ( .A1(n1690), .A2(n1691), .A3(n1692), .ZN(n1572) );
  NAND3_X1 U1343 ( .A1(n1690), .A2(n1691), .A3(n1692), .ZN(n1573) );
  XOR2_X1 U1344 ( .A(n367), .B(n380), .Z(n1574) );
  XOR2_X1 U1345 ( .A(n1489), .B(n1574), .Z(product[25]) );
  NAND2_X1 U1346 ( .A1(n1491), .A2(n367), .ZN(n1575) );
  NAND2_X1 U1347 ( .A1(n148), .A2(n380), .ZN(n1576) );
  NAND2_X1 U1348 ( .A1(n367), .A2(n380), .ZN(n1577) );
  NAND3_X1 U1349 ( .A1(n1575), .A2(n1576), .A3(n1577), .ZN(n147) );
  AND2_X1 U1350 ( .A1(n1829), .A2(b[16]), .ZN(n1578) );
  AND2_X1 U1351 ( .A1(n1832), .A2(b[15]), .ZN(n1579) );
  NOR3_X1 U1352 ( .A1(n1578), .A2(n1579), .A3(n2281), .ZN(n2280) );
  NAND2_X1 U1353 ( .A1(n1637), .A2(n2275), .ZN(n1580) );
  NAND2_X1 U1354 ( .A1(n1637), .A2(n473), .ZN(n1581) );
  NAND2_X1 U1355 ( .A1(n473), .A2(n2275), .ZN(n1582) );
  XOR2_X1 U1356 ( .A(n262), .B(n272), .Z(n1583) );
  XOR2_X1 U1357 ( .A(n1520), .B(n1583), .Z(product[33]) );
  NAND2_X1 U1358 ( .A1(n1542), .A2(n262), .ZN(n1584) );
  NAND2_X1 U1359 ( .A1(n140), .A2(n272), .ZN(n1585) );
  NAND2_X1 U1360 ( .A1(n262), .A2(n272), .ZN(n1586) );
  NAND3_X1 U1361 ( .A1(n1584), .A2(n1585), .A3(n1586), .ZN(n139) );
  CLKBUF_X1 U1362 ( .A(n649), .Z(n1587) );
  XOR2_X1 U1363 ( .A(n232), .B(n240), .Z(n1589) );
  XOR2_X1 U1364 ( .A(n1522), .B(n1589), .Z(product[36]) );
  NAND2_X1 U1365 ( .A1(n1543), .A2(n232), .ZN(n1590) );
  NAND2_X1 U1366 ( .A1(n137), .A2(n240), .ZN(n1591) );
  NAND2_X1 U1367 ( .A1(n232), .A2(n240), .ZN(n1592) );
  NAND3_X1 U1368 ( .A1(n1590), .A2(n1591), .A3(n1592), .ZN(n136) );
  XOR2_X1 U1369 ( .A(n485), .B(n860), .Z(n1593) );
  NAND2_X1 U1370 ( .A1(n492), .A2(n485), .ZN(n1594) );
  NAND2_X1 U1371 ( .A1(n492), .A2(n860), .ZN(n1595) );
  NAND2_X1 U1372 ( .A1(n485), .A2(n860), .ZN(n1596) );
  NAND3_X1 U1373 ( .A1(n1594), .A2(n1595), .A3(n1596), .ZN(n482) );
  XOR2_X1 U1374 ( .A(n846), .B(a[8]), .Z(n555) );
  NAND3_X1 U1375 ( .A1(n1653), .A2(n1654), .A3(n1655), .ZN(n1597) );
  NAND3_X1 U1376 ( .A1(n1653), .A2(n1654), .A3(n1655), .ZN(n1598) );
  NAND3_X1 U1377 ( .A1(n1693), .A2(n1694), .A3(n1695), .ZN(n1599) );
  OAI221_X1 U1378 ( .B1(n1841), .B2(n1947), .C1(n1837), .C2(n1784), .A(n1989), 
        .ZN(n1988) );
  NAND3_X2 U1379 ( .A1(n1488), .A2(n1993), .A3(n1996), .ZN(n1947) );
  INV_X1 U1380 ( .A(n665), .ZN(n1600) );
  CLKBUF_X1 U1381 ( .A(n1534), .Z(n1602) );
  CLKBUF_X1 U1382 ( .A(n135), .Z(n1603) );
  CLKBUF_X1 U1383 ( .A(n145), .Z(n1604) );
  XNOR2_X1 U1384 ( .A(n1605), .B(n174), .ZN(n1878) );
  NAND3_X1 U1385 ( .A1(n1748), .A2(n1747), .A3(n1749), .ZN(n1605) );
  INV_X1 U1386 ( .A(n1623), .ZN(n1789) );
  NAND2_X1 U1387 ( .A1(n1611), .A2(n1612), .ZN(n1993) );
  NAND2_X1 U1388 ( .A1(n2267), .A2(n2268), .ZN(n1606) );
  NAND2_X1 U1389 ( .A1(n2267), .A2(n449), .ZN(n1607) );
  NAND2_X1 U1390 ( .A1(n449), .A2(n2268), .ZN(n1608) );
  BUF_X4 U1391 ( .A(n1820), .Z(n1768) );
  BUF_X2 U1392 ( .A(n1814), .Z(n1766) );
  BUF_X2 U1393 ( .A(n1809), .Z(n1764) );
  BUF_X4 U1394 ( .A(n1825), .Z(n1771) );
  INV_X2 U1395 ( .A(n1884), .ZN(n1832) );
  XOR2_X1 U1396 ( .A(n532), .B(n1689), .Z(n527) );
  XOR2_X1 U1397 ( .A(n1515), .B(n1660), .Z(n676) );
  XOR2_X1 U1398 ( .A(n1601), .B(n1656), .Z(n680) );
  OR2_X1 U1399 ( .A1(a[7]), .A2(n1770), .ZN(n1612) );
  NAND3_X1 U1400 ( .A1(n1756), .A2(n1757), .A3(n1758), .ZN(n1609) );
  NAND3_X1 U1401 ( .A1(n1756), .A2(n1757), .A3(n1758), .ZN(n1610) );
  NAND2_X1 U1402 ( .A1(a[7]), .A2(n1770), .ZN(n1611) );
  BUF_X4 U1403 ( .A(n1825), .Z(n1770) );
  INV_X1 U1404 ( .A(n2246), .ZN(n1797) );
  INV_X1 U1405 ( .A(n2294), .ZN(n1830) );
  INV_X1 U1406 ( .A(n1473), .ZN(n1780) );
  INV_X1 U1407 ( .A(n1473), .ZN(n1781) );
  INV_X1 U1408 ( .A(n2218), .ZN(n1835) );
  INV_X1 U1409 ( .A(n2004), .ZN(n1819) );
  INV_X1 U1410 ( .A(n2171), .ZN(n1803) );
  INV_X1 U1411 ( .A(n2059), .ZN(n1813) );
  INV_X1 U1412 ( .A(n2115), .ZN(n1808) );
  INV_X1 U1413 ( .A(n2172), .ZN(n1805) );
  INV_X1 U1414 ( .A(n2060), .ZN(n1815) );
  INV_X1 U1415 ( .A(n2116), .ZN(n1810) );
  CLKBUF_X1 U1416 ( .A(n1944), .Z(n1784) );
  CLKBUF_X1 U1417 ( .A(n1999), .Z(n1788) );
  INV_X1 U1418 ( .A(n2002), .ZN(n1818) );
  INV_X1 U1419 ( .A(n2057), .ZN(n1812) );
  INV_X1 U1420 ( .A(n1947), .ZN(n1824) );
  INV_X1 U1421 ( .A(n2113), .ZN(n1807) );
  INV_X1 U1422 ( .A(n2169), .ZN(n1802) );
  NAND3_X1 U1423 ( .A1(n2217), .A2(n2216), .A3(n2221), .ZN(n2169) );
  NOR2_X2 U1424 ( .A1(n1811), .A2(n2164), .ZN(n2116) );
  NOR2_X2 U1425 ( .A1(n2160), .A2(n2161), .ZN(n2115) );
  INV_X1 U1426 ( .A(n2252), .ZN(n1795) );
  INV_X1 U1427 ( .A(n559), .ZN(n1826) );
  INV_X1 U1428 ( .A(n2223), .ZN(n1799) );
  INV_X1 U1429 ( .A(n545), .ZN(n1822) );
  INV_X1 U1430 ( .A(n533), .ZN(n1817) );
  INV_X1 U1431 ( .A(n553), .ZN(n1823) );
  INV_X1 U1432 ( .A(n1874), .ZN(n1649) );
  BUF_X1 U1433 ( .A(n1877), .Z(n1774) );
  BUF_X1 U1434 ( .A(n1877), .Z(n1775) );
  BUF_X1 U1435 ( .A(n2224), .Z(n1793) );
  BUF_X1 U1436 ( .A(n2224), .Z(n1794) );
  INV_X1 U1437 ( .A(n1888), .ZN(n1836) );
  BUF_X1 U1438 ( .A(n1804), .Z(n1762) );
  XNOR2_X1 U1439 ( .A(n436), .B(n1613), .ZN(n423) );
  XNOR2_X1 U1440 ( .A(n425), .B(n855), .ZN(n1613) );
  XNOR2_X1 U1441 ( .A(n1598), .B(n1614), .ZN(n449) );
  XNOR2_X1 U1442 ( .A(n451), .B(n857), .ZN(n1614) );
  XNOR2_X1 U1443 ( .A(n1569), .B(n1615), .ZN(n473) );
  XNOR2_X1 U1444 ( .A(n475), .B(n859), .ZN(n1615) );
  XNOR2_X1 U1445 ( .A(n544), .B(n1616), .ZN(n539) );
  XNOR2_X1 U1446 ( .A(n541), .B(n867), .ZN(n1616) );
  BUF_X2 U1447 ( .A(n1828), .Z(n1772) );
  BUF_X1 U1448 ( .A(n1820), .Z(n1769) );
  XNOR2_X1 U1449 ( .A(n463), .B(n858), .ZN(n1617) );
  BUF_X1 U1450 ( .A(n1809), .Z(n1765) );
  BUF_X1 U1451 ( .A(n1814), .Z(n1767) );
  BUF_X1 U1452 ( .A(n1804), .Z(n1763) );
  XNOR2_X1 U1453 ( .A(n521), .B(n864), .ZN(n1618) );
  XNOR2_X1 U1454 ( .A(n1599), .B(n1619), .ZN(n511) );
  XNOR2_X1 U1455 ( .A(n513), .B(n863), .ZN(n1619) );
  OAI221_X1 U1456 ( .B1(n1841), .B2(n2002), .C1(n1837), .C2(n1786), .A(n2044), 
        .ZN(n2043) );
  INV_X1 U1457 ( .A(n671), .ZN(n1846) );
  INV_X1 U1458 ( .A(n669), .ZN(n1843) );
  INV_X1 U1459 ( .A(n673), .ZN(n1849) );
  INV_X1 U1460 ( .A(n674), .ZN(n1851) );
  INV_X1 U1461 ( .A(n2217), .ZN(n1806) );
  INV_X1 U1462 ( .A(n2105), .ZN(n1816) );
  INV_X1 U1463 ( .A(n2161), .ZN(n1811) );
  INV_X1 U1464 ( .A(n684), .ZN(n1871) );
  INV_X1 U1465 ( .A(n682), .ZN(n1867) );
  INV_X1 U1466 ( .A(n675), .ZN(n1853) );
  INV_X1 U1467 ( .A(n685), .ZN(n1873) );
  INV_X1 U1468 ( .A(n677), .ZN(n1857) );
  INV_X1 U1469 ( .A(n679), .ZN(n1861) );
  INV_X1 U1470 ( .A(n681), .ZN(n1865) );
  INV_X1 U1471 ( .A(n676), .ZN(n1855) );
  INV_X1 U1472 ( .A(n680), .ZN(n1863) );
  INV_X1 U1473 ( .A(n683), .ZN(n1869) );
  INV_X1 U1474 ( .A(n678), .ZN(n1859) );
  INV_X1 U1475 ( .A(n434), .ZN(n1798) );
  INV_X1 U1476 ( .A(n686), .ZN(n1875) );
  INV_X1 U1477 ( .A(n2049), .ZN(n1821) );
  AND2_X1 U1478 ( .A1(n1806), .A2(n2216), .ZN(n1620) );
  AND2_X1 U1479 ( .A1(n1811), .A2(n2160), .ZN(n1621) );
  OR2_X1 U1480 ( .A1(n1821), .A2(n2052), .ZN(n1623) );
  INV_X1 U1481 ( .A(n2253), .ZN(n1800) );
  INV_X1 U1482 ( .A(n1893), .ZN(n1827) );
  INV_X1 U1483 ( .A(n1733), .ZN(n1881) );
  CLKBUF_X1 U1484 ( .A(n1890), .Z(n1779) );
  XOR2_X1 U1485 ( .A(a[4]), .B(n1828), .Z(n1624) );
  XOR2_X1 U1486 ( .A(a[3]), .B(a[2]), .Z(n1625) );
  INV_X1 U1487 ( .A(a[1]), .ZN(n1833) );
  INV_X1 U1488 ( .A(b[15]), .ZN(n1848) );
  INV_X1 U1489 ( .A(b[9]), .ZN(n1860) );
  INV_X1 U1490 ( .A(b[7]), .ZN(n1864) );
  INV_X1 U1491 ( .A(b[6]), .ZN(n1866) );
  INV_X1 U1492 ( .A(b[13]), .ZN(n1852) );
  INV_X1 U1493 ( .A(b[12]), .ZN(n1854) );
  INV_X1 U1494 ( .A(b[11]), .ZN(n1856) );
  INV_X1 U1495 ( .A(b[4]), .ZN(n1870) );
  INV_X1 U1496 ( .A(b[3]), .ZN(n1872) );
  INV_X1 U1497 ( .A(b[8]), .ZN(n1862) );
  INV_X1 U1498 ( .A(b[10]), .ZN(n1858) );
  INV_X1 U1499 ( .A(b[16]), .ZN(n1847) );
  INV_X1 U1500 ( .A(b[14]), .ZN(n1850) );
  INV_X1 U1501 ( .A(b[5]), .ZN(n1868) );
  XNOR2_X1 U1502 ( .A(n1513), .B(n1626), .ZN(n683) );
  XNOR2_X1 U1503 ( .A(b[3]), .B(b[4]), .ZN(n1626) );
  XNOR2_X1 U1504 ( .A(n1533), .B(n1627), .ZN(n678) );
  XNOR2_X1 U1505 ( .A(b[9]), .B(b[8]), .ZN(n1627) );
  NAND2_X1 U1506 ( .A1(a[1]), .A2(n1834), .ZN(n1884) );
  INV_X1 U1507 ( .A(b[2]), .ZN(n1874) );
  XOR2_X1 U1508 ( .A(n643), .B(n1629), .Z(n1628) );
  XNOR2_X1 U1509 ( .A(b[21]), .B(b[20]), .ZN(n1629) );
  XOR2_X1 U1510 ( .A(n1487), .B(n1631), .Z(n1630) );
  XNOR2_X1 U1511 ( .A(b[18]), .B(b[19]), .ZN(n1631) );
  XNOR2_X1 U1512 ( .A(b[14]), .B(b[15]), .ZN(n1633) );
  OAI221_X1 U1513 ( .B1(n1848), .B2(n2002), .C1(n1634), .C2(n1786), .A(n2034), 
        .ZN(n2033) );
  AOI221_X1 U1514 ( .B1(n1794), .B2(b[3]), .C1(n1797), .C2(n1649), .A(n2226), 
        .ZN(n709) );
  OAI221_X1 U1515 ( .B1(n1848), .B2(n2057), .C1(n1634), .C2(n1790), .A(n2090), 
        .ZN(n2089) );
  INV_X1 U1516 ( .A(a[17]), .ZN(n1809) );
  INV_X1 U1517 ( .A(a[20]), .ZN(n1804) );
  INV_X1 U1518 ( .A(a[14]), .ZN(n1814) );
  INV_X1 U1519 ( .A(a[0]), .ZN(n1834) );
  INV_X1 U1520 ( .A(a[11]), .ZN(n1820) );
  INV_X1 U1521 ( .A(a[8]), .ZN(n1825) );
  INV_X1 U1522 ( .A(b[0]), .ZN(n1877) );
  OAI221_X1 U1523 ( .B1(n1848), .B2(n2169), .C1(n1634), .C2(n1792), .A(n2202), 
        .ZN(n2201) );
  OAI221_X1 U1524 ( .B1(n1848), .B2(n2113), .C1(n1634), .C2(n1791), .A(n2146), 
        .ZN(n2145) );
  INV_X1 U1525 ( .A(b[19]), .ZN(n1842) );
  INV_X1 U1526 ( .A(b[18]), .ZN(n1844) );
  INV_X1 U1527 ( .A(b[17]), .ZN(n1845) );
  INV_X1 U1528 ( .A(b[20]), .ZN(n1841) );
  INV_X1 U1529 ( .A(b[22]), .ZN(n1838) );
  NAND2_X1 U1530 ( .A1(n1829), .A2(b[22]), .ZN(n1635) );
  NAND2_X1 U1531 ( .A1(n1832), .A2(b[21]), .ZN(n1636) );
  INV_X1 U1532 ( .A(b[21]), .ZN(n1839) );
  XNOR2_X1 U1533 ( .A(n1878), .B(n1839), .ZN(product[47]) );
  OAI222_X1 U1534 ( .A1(n2279), .A2(n2278), .B1(n2278), .B2(n1477), .C1(n2279), 
        .C2(n1477), .ZN(n1637) );
  NAND2_X1 U1535 ( .A1(n2290), .A2(n2291), .ZN(n1638) );
  NAND2_X1 U1536 ( .A1(n2290), .A2(n511), .ZN(n1639) );
  NAND2_X1 U1537 ( .A1(n511), .A2(n2291), .ZN(n1640) );
  NAND2_X1 U1538 ( .A1(n1599), .A2(n513), .ZN(n1641) );
  NAND2_X1 U1539 ( .A1(n518), .A2(n863), .ZN(n1642) );
  NAND2_X1 U1540 ( .A1(n513), .A2(n863), .ZN(n1643) );
  NAND3_X1 U1541 ( .A1(n1641), .A2(n1642), .A3(n1643), .ZN(n510) );
  NAND2_X1 U1542 ( .A1(n1597), .A2(n451), .ZN(n1644) );
  NAND2_X1 U1543 ( .A1(n460), .A2(n857), .ZN(n1645) );
  NAND2_X1 U1544 ( .A1(n451), .A2(n857), .ZN(n1646) );
  NAND3_X1 U1545 ( .A1(n1644), .A2(n1645), .A3(n1646), .ZN(n448) );
  XNOR2_X1 U1546 ( .A(a[3]), .B(a[2]), .ZN(n1647) );
  NAND2_X1 U1547 ( .A1(n436), .A2(n425), .ZN(n1650) );
  NAND2_X1 U1548 ( .A1(n436), .A2(n855), .ZN(n1651) );
  NAND2_X1 U1549 ( .A1(n425), .A2(n855), .ZN(n1652) );
  NAND3_X1 U1550 ( .A1(n1651), .A2(n1650), .A3(n1652), .ZN(n422) );
  NAND2_X1 U1551 ( .A1(n1570), .A2(n463), .ZN(n1653) );
  NAND2_X1 U1552 ( .A1(n472), .A2(n858), .ZN(n1654) );
  NAND2_X1 U1553 ( .A1(n463), .A2(n858), .ZN(n1655) );
  NAND3_X1 U1554 ( .A1(n1653), .A2(n1654), .A3(n1655), .ZN(n460) );
  XOR2_X1 U1555 ( .A(b[0]), .B(n1519), .Z(n686) );
  XOR2_X1 U1556 ( .A(b[7]), .B(b[6]), .Z(n1656) );
  NAND2_X1 U1557 ( .A1(n657), .A2(b[7]), .ZN(n1657) );
  NAND2_X1 U1558 ( .A1(n657), .A2(b[6]), .ZN(n1658) );
  NAND2_X1 U1559 ( .A1(b[7]), .A2(b[6]), .ZN(n1659) );
  NAND3_X1 U1560 ( .A1(n1657), .A2(n1658), .A3(n1659), .ZN(n656) );
  XOR2_X1 U1561 ( .A(b[10]), .B(b[11]), .Z(n1660) );
  NAND2_X1 U1562 ( .A1(n653), .A2(b[10]), .ZN(n1661) );
  NAND2_X1 U1563 ( .A1(n653), .A2(b[11]), .ZN(n1662) );
  NAND2_X1 U1564 ( .A1(b[10]), .A2(b[11]), .ZN(n1663) );
  NAND3_X1 U1565 ( .A1(n1661), .A2(n1662), .A3(n1663), .ZN(n652) );
  NAND2_X1 U1566 ( .A1(n660), .A2(b[3]), .ZN(n1664) );
  NAND2_X1 U1567 ( .A1(n660), .A2(b[4]), .ZN(n1665) );
  NAND2_X1 U1568 ( .A1(b[3]), .A2(b[4]), .ZN(n1666) );
  NAND3_X1 U1569 ( .A1(n1665), .A2(n1664), .A3(n1666), .ZN(n659) );
  XOR2_X1 U1570 ( .A(b[16]), .B(b[17]), .Z(n1667) );
  NAND2_X1 U1571 ( .A1(n647), .A2(b[16]), .ZN(n1668) );
  NAND2_X1 U1572 ( .A1(n647), .A2(b[17]), .ZN(n1669) );
  NAND2_X1 U1573 ( .A1(b[16]), .A2(b[17]), .ZN(n1670) );
  NAND3_X1 U1574 ( .A1(n1669), .A2(n1668), .A3(n1670), .ZN(n646) );
  NAND2_X1 U1575 ( .A1(n643), .A2(b[21]), .ZN(n1671) );
  NAND2_X1 U1576 ( .A1(n643), .A2(b[20]), .ZN(n1672) );
  NAND2_X1 U1577 ( .A1(b[21]), .A2(b[20]), .ZN(n1673) );
  NAND3_X1 U1578 ( .A1(n1671), .A2(n1672), .A3(n1673), .ZN(n642) );
  AND2_X1 U1579 ( .A1(n1829), .A2(b[18]), .ZN(n1674) );
  AND2_X1 U1580 ( .A1(n1832), .A2(b[17]), .ZN(n1675) );
  NOR3_X1 U1581 ( .A1(n1674), .A2(n1675), .A3(n2274), .ZN(n2273) );
  NAND2_X1 U1582 ( .A1(n2282), .A2(n2283), .ZN(n1676) );
  NAND2_X1 U1583 ( .A1(n2282), .A2(n493), .ZN(n1677) );
  NAND2_X1 U1584 ( .A1(n493), .A2(n2283), .ZN(n1678) );
  NAND2_X1 U1585 ( .A1(n2315), .A2(n2316), .ZN(n1679) );
  NAND2_X1 U1586 ( .A1(n2315), .A2(n549), .ZN(n1680) );
  NAND2_X1 U1587 ( .A1(n549), .A2(n2316), .ZN(n1681) );
  INV_X1 U1588 ( .A(n1534), .ZN(n1876) );
  AND3_X1 U1589 ( .A1(n1718), .A2(n1717), .A3(n1719), .ZN(n1682) );
  AND2_X1 U1590 ( .A1(n1829), .A2(b[17]), .ZN(n1683) );
  AND2_X1 U1591 ( .A1(n1832), .A2(b[16]), .ZN(n1684) );
  NOR3_X1 U1592 ( .A1(n1683), .A2(n1684), .A3(n2277), .ZN(n2276) );
  XOR2_X1 U1593 ( .A(n325), .B(n338), .Z(n1685) );
  XOR2_X1 U1594 ( .A(n1604), .B(n1685), .Z(product[28]) );
  NAND2_X1 U1595 ( .A1(n145), .A2(n325), .ZN(n1686) );
  NAND2_X1 U1596 ( .A1(n1523), .A2(n338), .ZN(n1687) );
  NAND2_X1 U1597 ( .A1(n325), .A2(n338), .ZN(n1688) );
  NAND3_X1 U1598 ( .A1(n1686), .A2(n1687), .A3(n1688), .ZN(n144) );
  XOR2_X1 U1599 ( .A(n529), .B(n865), .Z(n1689) );
  NAND2_X1 U1600 ( .A1(n532), .A2(n529), .ZN(n1690) );
  NAND2_X1 U1601 ( .A1(n532), .A2(n865), .ZN(n1691) );
  NAND2_X1 U1602 ( .A1(n529), .A2(n865), .ZN(n1692) );
  NAND3_X1 U1603 ( .A1(n1690), .A2(n1691), .A3(n1692), .ZN(n526) );
  NAND2_X1 U1604 ( .A1(n1572), .A2(n521), .ZN(n1693) );
  NAND2_X1 U1605 ( .A1(n526), .A2(n864), .ZN(n1694) );
  NAND2_X1 U1606 ( .A1(n521), .A2(n864), .ZN(n1695) );
  NAND3_X1 U1607 ( .A1(n1693), .A2(n1694), .A3(n1695), .ZN(n518) );
  XOR2_X1 U1608 ( .A(n284), .B(n273), .Z(n1696) );
  XOR2_X1 U1609 ( .A(n1610), .B(n1696), .Z(product[32]) );
  NAND2_X1 U1610 ( .A1(n1609), .A2(n284), .ZN(n1697) );
  NAND2_X1 U1611 ( .A1(n141), .A2(n273), .ZN(n1698) );
  NAND2_X1 U1612 ( .A1(n284), .A2(n273), .ZN(n1699) );
  NAND3_X1 U1613 ( .A1(n1698), .A2(n1697), .A3(n1699), .ZN(n140) );
  AND2_X1 U1614 ( .A1(n1829), .A2(b[20]), .ZN(n1700) );
  AND2_X1 U1615 ( .A1(n1832), .A2(b[19]), .ZN(n1701) );
  INV_X1 U1616 ( .A(n437), .ZN(n1801) );
  NAND2_X1 U1617 ( .A1(n649), .A2(b[14]), .ZN(n1702) );
  NAND2_X1 U1618 ( .A1(n649), .A2(b[15]), .ZN(n1703) );
  NAND2_X1 U1619 ( .A1(b[14]), .A2(b[15]), .ZN(n1704) );
  NAND3_X1 U1620 ( .A1(n1702), .A2(n1703), .A3(n1704), .ZN(n648) );
  CLKBUF_X1 U1621 ( .A(n138), .Z(n1705) );
  AND2_X1 U1622 ( .A1(n1829), .A2(b[21]), .ZN(n1706) );
  AND2_X1 U1623 ( .A1(n1832), .A2(b[20]), .ZN(n1707) );
  NOR3_X1 U1624 ( .A1(n1706), .A2(n1707), .A3(n2262), .ZN(n2261) );
  XNOR2_X1 U1625 ( .A(n1918), .B(n1772), .ZN(n859) );
  INV_X1 U1626 ( .A(a[5]), .ZN(n1828) );
  XOR2_X1 U1627 ( .A(n250), .B(n241), .Z(n1708) );
  XOR2_X1 U1628 ( .A(n1705), .B(n1708), .Z(product[35]) );
  NAND2_X1 U1629 ( .A1(n138), .A2(n250), .ZN(n1709) );
  NAND2_X1 U1630 ( .A1(n138), .A2(n241), .ZN(n1710) );
  NAND2_X1 U1631 ( .A1(n250), .A2(n241), .ZN(n1711) );
  NAND3_X1 U1632 ( .A1(n1710), .A2(n1709), .A3(n1711), .ZN(n137) );
  NOR2_X1 U1633 ( .A1(n2258), .A2(n1480), .ZN(n2257) );
  INV_X1 U1634 ( .A(n665), .ZN(n1837) );
  XOR2_X1 U1635 ( .A(n222), .B(n215), .Z(n1712) );
  XOR2_X1 U1636 ( .A(n1603), .B(n1712), .Z(product[38]) );
  NAND2_X1 U1637 ( .A1(n135), .A2(n222), .ZN(n1713) );
  NAND2_X1 U1638 ( .A1(n135), .A2(n215), .ZN(n1714) );
  NAND2_X1 U1639 ( .A1(n222), .A2(n215), .ZN(n1715) );
  NAND3_X1 U1640 ( .A1(n1713), .A2(n1714), .A3(n1715), .ZN(n134) );
  INV_X1 U1641 ( .A(n1776), .ZN(n1716) );
  NAND2_X1 U1642 ( .A1(n2259), .A2(n2260), .ZN(n1717) );
  NAND2_X1 U1643 ( .A1(n2259), .A2(n423), .ZN(n1718) );
  NAND2_X1 U1644 ( .A1(n2260), .A2(n423), .ZN(n1719) );
  AND3_X1 U1645 ( .A1(n1717), .A2(n1718), .A3(n1719), .ZN(n2255) );
  CLKBUF_X1 U1646 ( .A(n1877), .Z(n1776) );
  XOR2_X1 U1647 ( .A(n201), .B(n207), .Z(n1720) );
  XOR2_X1 U1648 ( .A(n1539), .B(n1720), .Z(product[40]) );
  NAND2_X1 U1649 ( .A1(n133), .A2(n201), .ZN(n1721) );
  NAND2_X1 U1650 ( .A1(n133), .A2(n207), .ZN(n1722) );
  NAND2_X1 U1651 ( .A1(n201), .A2(n207), .ZN(n1723) );
  NAND3_X1 U1652 ( .A1(n1722), .A2(n1721), .A3(n1723), .ZN(n132) );
  XOR2_X1 U1653 ( .A(n381), .B(n876), .Z(n1724) );
  XOR2_X1 U1654 ( .A(n1521), .B(n1724), .Z(product[24]) );
  NAND2_X1 U1655 ( .A1(n149), .A2(n381), .ZN(n1725) );
  NAND2_X1 U1656 ( .A1(n149), .A2(n876), .ZN(n1726) );
  NAND2_X1 U1657 ( .A1(n381), .A2(n876), .ZN(n1727) );
  NAND3_X1 U1658 ( .A1(n1726), .A2(n1725), .A3(n1727), .ZN(n148) );
  NAND2_X1 U1659 ( .A1(n544), .A2(n541), .ZN(n1728) );
  NAND2_X1 U1660 ( .A1(n544), .A2(n867), .ZN(n1729) );
  NAND2_X1 U1661 ( .A1(n541), .A2(n867), .ZN(n1730) );
  NAND3_X1 U1662 ( .A1(n1728), .A2(n1729), .A3(n1730), .ZN(n538) );
  XNOR2_X1 U1663 ( .A(a[4]), .B(n1828), .ZN(n1731) );
  XNOR2_X1 U1664 ( .A(a[4]), .B(n1773), .ZN(n1732) );
  OR3_X4 U1665 ( .A1(n2335), .A2(a[0]), .A3(a[1]), .ZN(n1733) );
  XOR2_X1 U1666 ( .A(n190), .B(n194), .Z(n1734) );
  XOR2_X1 U1667 ( .A(n1738), .B(n1734), .Z(product[42]) );
  NAND2_X1 U1668 ( .A1(n131), .A2(n190), .ZN(n1735) );
  NAND2_X1 U1669 ( .A1(n131), .A2(n194), .ZN(n1736) );
  NAND2_X1 U1670 ( .A1(n190), .A2(n194), .ZN(n1737) );
  NAND3_X1 U1671 ( .A1(n1736), .A2(n1735), .A3(n1737), .ZN(n130) );
  CLKBUF_X1 U1672 ( .A(n131), .Z(n1738) );
  NAND2_X1 U1673 ( .A1(n645), .A2(b[18]), .ZN(n1739) );
  NAND2_X1 U1674 ( .A1(n645), .A2(b[19]), .ZN(n1740) );
  NAND2_X1 U1675 ( .A1(b[18]), .A2(b[19]), .ZN(n1741) );
  NAND3_X1 U1676 ( .A1(n1740), .A2(n1739), .A3(n1741), .ZN(n644) );
  NAND2_X1 U1677 ( .A1(n655), .A2(b[9]), .ZN(n1742) );
  NAND2_X1 U1678 ( .A1(n655), .A2(b[8]), .ZN(n1743) );
  NAND2_X1 U1679 ( .A1(b[9]), .A2(b[8]), .ZN(n1744) );
  NAND3_X1 U1680 ( .A1(n1743), .A2(n1742), .A3(n1744), .ZN(n654) );
  CLKBUF_X1 U1681 ( .A(n1602), .Z(n1745) );
  INV_X1 U1682 ( .A(n409), .ZN(n1796) );
  XOR2_X1 U1683 ( .A(n175), .B(n177), .Z(n1746) );
  XOR2_X1 U1684 ( .A(n1750), .B(n1746), .Z(product[46]) );
  NAND2_X1 U1685 ( .A1(n127), .A2(n175), .ZN(n1747) );
  NAND2_X1 U1686 ( .A1(n127), .A2(n177), .ZN(n1748) );
  NAND2_X1 U1687 ( .A1(n175), .A2(n177), .ZN(n1749) );
  CLKBUF_X1 U1688 ( .A(n127), .Z(n1750) );
  XOR2_X1 U1689 ( .A(n184), .B(n181), .Z(n1751) );
  XOR2_X1 U1690 ( .A(n1540), .B(n1751), .Z(product[44]) );
  NAND2_X1 U1691 ( .A1(n129), .A2(n184), .ZN(n1752) );
  NAND2_X1 U1692 ( .A1(n129), .A2(n181), .ZN(n1753) );
  NAND2_X1 U1693 ( .A1(n184), .A2(n181), .ZN(n1754) );
  NAND3_X1 U1694 ( .A1(n1752), .A2(n1753), .A3(n1754), .ZN(n128) );
  XOR2_X1 U1695 ( .A(n285), .B(n297), .Z(n1755) );
  XOR2_X1 U1696 ( .A(n1541), .B(n1755), .Z(product[31]) );
  NAND2_X1 U1697 ( .A1(n142), .A2(n285), .ZN(n1756) );
  NAND2_X1 U1698 ( .A1(n142), .A2(n297), .ZN(n1757) );
  NAND2_X1 U1699 ( .A1(n285), .A2(n297), .ZN(n1758) );
  NAND3_X1 U1700 ( .A1(n1756), .A2(n1757), .A3(n1758), .ZN(n141) );
  NAND2_X1 U1701 ( .A1(n1568), .A2(n475), .ZN(n1759) );
  NAND2_X1 U1702 ( .A1(n482), .A2(n859), .ZN(n1760) );
  NAND2_X1 U1703 ( .A1(n475), .A2(n859), .ZN(n1761) );
  NAND3_X1 U1704 ( .A1(n1759), .A2(n1760), .A3(n1761), .ZN(n472) );
  BUF_X4 U1705 ( .A(n1828), .Z(n1773) );
  BUF_X2 U1706 ( .A(n1890), .Z(n1778) );
  BUF_X2 U1707 ( .A(n1999), .Z(n1786) );
  BUF_X2 U1708 ( .A(n1999), .Z(n1787) );
  NOR2_X4 U1709 ( .A1(n2048), .A2(n2049), .ZN(n2004) );
  NAND3_X2 U1710 ( .A1(n2049), .A2(n2048), .A3(n2052), .ZN(n2002) );
  NOR2_X4 U1711 ( .A1(n2104), .A2(n2105), .ZN(n2059) );
  NOR2_X4 U1712 ( .A1(n1816), .A2(n2108), .ZN(n2060) );
  NAND3_X2 U1713 ( .A1(n2105), .A2(n2104), .A3(n2108), .ZN(n2057) );
  NAND3_X2 U1714 ( .A1(n2161), .A2(n2160), .A3(n2164), .ZN(n2113) );
  NOR2_X4 U1715 ( .A1(n2216), .A2(n2217), .ZN(n2171) );
  NOR2_X4 U1716 ( .A1(n1806), .A2(n2221), .ZN(n2172) );
  INV_X1 U1717 ( .A(n1472), .ZN(n1790) );
  INV_X1 U1718 ( .A(n1621), .ZN(n1791) );
  INV_X1 U1719 ( .A(n1620), .ZN(n1792) );
  XNOR2_X1 U1720 ( .A(n1879), .B(n1496), .ZN(n877) );
  OAI21_X1 U1721 ( .B1(n1492), .B2(n1830), .A(n1880), .ZN(n1879) );
  OAI22_X1 U1722 ( .A1(n1881), .A2(n1882), .B1(b[21]), .B2(n1882), .ZN(n1880)
         );
  AOI22_X1 U1723 ( .A1(n1883), .A2(n1884), .B1(n1883), .B2(n1838), .ZN(n1882)
         );
  XNOR2_X1 U1724 ( .A(n1885), .B(n1496), .ZN(n876) );
  OAI21_X1 U1725 ( .B1(n1830), .B2(n1836), .A(n1886), .ZN(n1885) );
  OAI22_X1 U1726 ( .A1(n1881), .A2(n1832), .B1(b[22]), .B2(n1832), .ZN(n1886)
         );
  XNOR2_X1 U1727 ( .A(n1887), .B(n1496), .ZN(n875) );
  OAI21_X1 U1728 ( .B1(n1888), .B2(n1830), .A(n1733), .ZN(n1887) );
  XNOR2_X1 U1729 ( .A(n1889), .B(n1772), .ZN(n873) );
  OAI22_X1 U1730 ( .A1(n1774), .A2(n1484), .B1(n1777), .B2(n1775), .ZN(n1889)
         );
  XNOR2_X1 U1731 ( .A(n1891), .B(n1773), .ZN(n872) );
  OAI222_X1 U1732 ( .A1(n1776), .A2(n1473), .B1(n1484), .B2(n1876), .C1(n1778), 
        .C2(n1875), .ZN(n1891) );
  XNOR2_X1 U1733 ( .A(n1892), .B(n1772), .ZN(n871) );
  OAI221_X1 U1734 ( .B1(n1774), .B2(n1893), .C1(n1778), .C2(n1873), .A(n1894), 
        .ZN(n1892) );
  AOI22_X1 U1735 ( .A1(b[2]), .A2(n1895), .B1(n1781), .B2(n1602), .ZN(n1894)
         );
  XNOR2_X1 U1736 ( .A(n1896), .B(n1773), .ZN(n870) );
  OAI221_X1 U1737 ( .B1(n1876), .B2(n1893), .C1(n1778), .C2(n1871), .A(n1897), 
        .ZN(n1896) );
  AOI22_X1 U1738 ( .A1(b[3]), .A2(n1895), .B1(n1649), .B2(n1780), .ZN(n1897)
         );
  XNOR2_X1 U1739 ( .A(n1898), .B(n1772), .ZN(n869) );
  OAI221_X1 U1740 ( .B1(n1874), .B2(n1893), .C1(n1778), .C2(n1869), .A(n1899), 
        .ZN(n1898) );
  AOI22_X1 U1741 ( .A1(b[4]), .A2(n1895), .B1(b[3]), .B2(n1780), .ZN(n1899) );
  XNOR2_X1 U1742 ( .A(n1900), .B(n1773), .ZN(n868) );
  OAI221_X1 U1743 ( .B1(n1893), .B2(n1872), .C1(n1778), .C2(n1867), .A(n1901), 
        .ZN(n1900) );
  AOI22_X1 U1744 ( .A1(b[5]), .A2(n1895), .B1(b[4]), .B2(n1780), .ZN(n1901) );
  XNOR2_X1 U1745 ( .A(n1902), .B(n1772), .ZN(n867) );
  OAI221_X1 U1746 ( .B1(n1893), .B2(n1870), .C1(n1778), .C2(n1865), .A(n1903), 
        .ZN(n1902) );
  AOI22_X1 U1747 ( .A1(n1895), .A2(b[6]), .B1(b[5]), .B2(n1780), .ZN(n1903) );
  XNOR2_X1 U1748 ( .A(n1904), .B(n1773), .ZN(n866) );
  OAI221_X1 U1749 ( .B1(n1483), .B2(n1868), .C1(n1778), .C2(n1863), .A(n1905), 
        .ZN(n1904) );
  AOI22_X1 U1750 ( .A1(n1895), .A2(b[7]), .B1(n1781), .B2(b[6]), .ZN(n1905) );
  XNOR2_X1 U1751 ( .A(n1906), .B(n1772), .ZN(n865) );
  OAI221_X1 U1752 ( .B1(n1866), .B2(n1483), .C1(n1778), .C2(n1861), .A(n1907), 
        .ZN(n1906) );
  AOI22_X1 U1753 ( .A1(b[8]), .A2(n1895), .B1(n1781), .B2(b[7]), .ZN(n1907) );
  XNOR2_X1 U1754 ( .A(n1908), .B(n1773), .ZN(n864) );
  OAI221_X1 U1755 ( .B1(n1864), .B2(n1483), .C1(n1778), .C2(n1859), .A(n1909), 
        .ZN(n1908) );
  AOI22_X1 U1756 ( .A1(n1895), .A2(b[9]), .B1(b[8]), .B2(n1780), .ZN(n1909) );
  XNOR2_X1 U1757 ( .A(n1910), .B(n1772), .ZN(n863) );
  OAI221_X1 U1758 ( .B1(n1483), .B2(n1862), .C1(n1778), .C2(n1857), .A(n1911), 
        .ZN(n1910) );
  AOI22_X1 U1759 ( .A1(b[10]), .A2(n1895), .B1(n1781), .B2(b[9]), .ZN(n1911)
         );
  OAI221_X1 U1760 ( .B1(n1860), .B2(n1483), .C1(n1778), .C2(n1855), .A(n1913), 
        .ZN(n1912) );
  AOI22_X1 U1761 ( .A1(b[11]), .A2(n1895), .B1(b[10]), .B2(n1780), .ZN(n1913)
         );
  XNOR2_X1 U1762 ( .A(n1914), .B(n1772), .ZN(n861) );
  OAI221_X1 U1763 ( .B1(n1483), .B2(n1858), .C1(n1777), .C2(n1853), .A(n1915), 
        .ZN(n1914) );
  AOI22_X1 U1764 ( .A1(n1895), .A2(b[12]), .B1(b[11]), .B2(n1780), .ZN(n1915)
         );
  XNOR2_X1 U1765 ( .A(n1916), .B(n1773), .ZN(n860) );
  OAI221_X1 U1766 ( .B1(n1483), .B2(n1856), .C1(n1777), .C2(n1851), .A(n1917), 
        .ZN(n1916) );
  AOI22_X1 U1767 ( .A1(n1895), .A2(b[13]), .B1(n1781), .B2(b[12]), .ZN(n1917)
         );
  OAI221_X1 U1768 ( .B1(n1854), .B2(n1483), .C1(n1777), .C2(n1849), .A(n1919), 
        .ZN(n1918) );
  AOI22_X1 U1769 ( .A1(b[14]), .A2(n1895), .B1(n1781), .B2(b[13]), .ZN(n1919)
         );
  XNOR2_X1 U1770 ( .A(n1920), .B(n1773), .ZN(n858) );
  AOI22_X1 U1771 ( .A1(n1895), .A2(b[15]), .B1(b[14]), .B2(n1780), .ZN(n1921)
         );
  XNOR2_X1 U1772 ( .A(n1922), .B(n1772), .ZN(n857) );
  OAI221_X1 U1773 ( .B1(n1483), .B2(n1850), .C1(n1777), .C2(n1846), .A(n1923), 
        .ZN(n1922) );
  AOI22_X1 U1774 ( .A1(b[16]), .A2(n1895), .B1(n1781), .B2(b[15]), .ZN(n1923)
         );
  XNOR2_X1 U1775 ( .A(n1924), .B(n1773), .ZN(n856) );
  AOI22_X1 U1776 ( .A1(b[17]), .A2(n1895), .B1(b[16]), .B2(n1780), .ZN(n1925)
         );
  XNOR2_X1 U1777 ( .A(n1926), .B(n1773), .ZN(n855) );
  OAI221_X1 U1778 ( .B1(n1483), .B2(n1847), .C1(n1777), .C2(n1843), .A(n1927), 
        .ZN(n1926) );
  AOI22_X1 U1779 ( .A1(n1895), .A2(b[18]), .B1(b[17]), .B2(n1780), .ZN(n1927)
         );
  XNOR2_X1 U1780 ( .A(n1928), .B(n1772), .ZN(n854) );
  OAI221_X1 U1781 ( .B1(n1483), .B2(n1845), .C1(n1777), .C2(n1630), .A(n1929), 
        .ZN(n1928) );
  AOI22_X1 U1782 ( .A1(n1895), .A2(b[19]), .B1(n1781), .B2(b[18]), .ZN(n1929)
         );
  XNOR2_X1 U1783 ( .A(n1930), .B(n1773), .ZN(n853) );
  OAI221_X1 U1784 ( .B1(n1844), .B2(n1483), .C1(n1777), .C2(n1840), .A(n1931), 
        .ZN(n1930) );
  AOI22_X1 U1785 ( .A1(b[20]), .A2(n1895), .B1(n1781), .B2(b[19]), .ZN(n1931)
         );
  XNOR2_X1 U1786 ( .A(n1932), .B(n1772), .ZN(n852) );
  OAI221_X1 U1787 ( .B1(n1842), .B2(n1483), .C1(n1777), .C2(n1628), .A(n1933), 
        .ZN(n1932) );
  AOI22_X1 U1788 ( .A1(n1895), .A2(b[21]), .B1(b[20]), .B2(n1780), .ZN(n1933)
         );
  XNOR2_X1 U1789 ( .A(n1934), .B(n1773), .ZN(n851) );
  OAI221_X1 U1790 ( .B1(n1483), .B2(n1841), .C1(n1777), .C2(n1837), .A(n1935), 
        .ZN(n1934) );
  AOI22_X1 U1791 ( .A1(n1895), .A2(b[22]), .B1(n1781), .B2(b[21]), .ZN(n1935)
         );
  XNOR2_X1 U1792 ( .A(n1936), .B(n1772), .ZN(n850) );
  OAI21_X1 U1793 ( .B1(n1835), .B2(n1778), .A(n1937), .ZN(n1936) );
  OAI22_X1 U1794 ( .A1(n1827), .A2(n1938), .B1(b[21]), .B2(n1938), .ZN(n1937)
         );
  AOI22_X1 U1795 ( .A1(n1473), .A2(n1484), .B1(n1838), .B2(n1484), .ZN(n1938)
         );
  XNOR2_X1 U1796 ( .A(n1939), .B(n1773), .ZN(n849) );
  OAI21_X1 U1797 ( .B1(n1836), .B2(n1779), .A(n1940), .ZN(n1939) );
  OAI22_X1 U1798 ( .A1(n1827), .A2(n1781), .B1(b[22]), .B2(n1780), .ZN(n1940)
         );
  XNOR2_X1 U1799 ( .A(n1942), .B(n1772), .ZN(n848) );
  OAI21_X1 U1800 ( .B1(n1888), .B2(n1779), .A(n1483), .ZN(n1942) );
  XNOR2_X1 U1801 ( .A(a[3]), .B(a[4]), .ZN(n1941) );
  NAND2_X1 U1802 ( .A1(n1625), .A2(n1731), .ZN(n1890) );
  XNOR2_X1 U1803 ( .A(n1943), .B(n1770), .ZN(n846) );
  OAI22_X1 U1804 ( .A1(n1774), .A2(n1588), .B1(n1775), .B2(n1782), .ZN(n1943)
         );
  XNOR2_X1 U1805 ( .A(n1945), .B(n1771), .ZN(n845) );
  OAI222_X1 U1806 ( .A1(n1775), .A2(n1622), .B1(n1876), .B2(n1588), .C1(n1875), 
        .C2(n1782), .ZN(n1945) );
  XNOR2_X1 U1807 ( .A(n1946), .B(n1771), .ZN(n844) );
  OAI221_X1 U1808 ( .B1(n1774), .B2(n1947), .C1(n1873), .C2(n1783), .A(n1948), 
        .ZN(n1946) );
  AOI22_X1 U1809 ( .A1(n1949), .A2(n1649), .B1(n1785), .B2(n1602), .ZN(n1948)
         );
  XNOR2_X1 U1810 ( .A(n1950), .B(n1771), .ZN(n843) );
  OAI221_X1 U1811 ( .B1(n1876), .B2(n1947), .C1(n1871), .C2(n1784), .A(n1951), 
        .ZN(n1950) );
  AOI22_X1 U1812 ( .A1(n1949), .A2(b[3]), .B1(n1785), .B2(n1649), .ZN(n1951)
         );
  XNOR2_X1 U1813 ( .A(n1952), .B(n1771), .ZN(n842) );
  OAI221_X1 U1814 ( .B1(n1874), .B2(n1947), .C1(n1869), .C2(n1783), .A(n1953), 
        .ZN(n1952) );
  AOI22_X1 U1815 ( .A1(n1949), .A2(b[4]), .B1(n1785), .B2(b[3]), .ZN(n1953) );
  XNOR2_X1 U1816 ( .A(n1954), .B(n1771), .ZN(n841) );
  OAI221_X1 U1817 ( .B1(n1872), .B2(n1947), .C1(n1867), .C2(n1783), .A(n1955), 
        .ZN(n1954) );
  AOI22_X1 U1818 ( .A1(n1949), .A2(b[5]), .B1(n1785), .B2(b[4]), .ZN(n1955) );
  XNOR2_X1 U1819 ( .A(n1956), .B(n1771), .ZN(n840) );
  OAI221_X1 U1820 ( .B1(n1870), .B2(n1947), .C1(n1865), .C2(n1784), .A(n1957), 
        .ZN(n1956) );
  AOI22_X1 U1821 ( .A1(n1949), .A2(b[6]), .B1(n1785), .B2(b[5]), .ZN(n1957) );
  XNOR2_X1 U1822 ( .A(n1958), .B(n1771), .ZN(n839) );
  OAI221_X1 U1823 ( .B1(n1868), .B2(n1947), .C1(n1863), .C2(n1783), .A(n1959), 
        .ZN(n1958) );
  AOI22_X1 U1824 ( .A1(n1949), .A2(b[7]), .B1(n1785), .B2(b[6]), .ZN(n1959) );
  XNOR2_X1 U1825 ( .A(n1960), .B(n1771), .ZN(n838) );
  OAI221_X1 U1826 ( .B1(n1866), .B2(n1947), .C1(n1861), .C2(n1784), .A(n1961), 
        .ZN(n1960) );
  AOI22_X1 U1827 ( .A1(n1949), .A2(b[8]), .B1(n1785), .B2(b[7]), .ZN(n1961) );
  XNOR2_X1 U1828 ( .A(n1962), .B(n1771), .ZN(n837) );
  OAI221_X1 U1829 ( .B1(n1864), .B2(n1947), .C1(n1859), .C2(n1783), .A(n1963), 
        .ZN(n1962) );
  AOI22_X1 U1830 ( .A1(n1949), .A2(b[9]), .B1(n1785), .B2(b[8]), .ZN(n1963) );
  XNOR2_X1 U1831 ( .A(n1964), .B(n1771), .ZN(n836) );
  OAI221_X1 U1832 ( .B1(n1862), .B2(n1947), .C1(n1857), .C2(n1783), .A(n1965), 
        .ZN(n1964) );
  AOI22_X1 U1833 ( .A1(n1949), .A2(b[10]), .B1(n1785), .B2(b[9]), .ZN(n1965)
         );
  XNOR2_X1 U1834 ( .A(n1966), .B(n1771), .ZN(n835) );
  OAI221_X1 U1835 ( .B1(n1860), .B2(n1947), .C1(n1855), .C2(n1783), .A(n1967), 
        .ZN(n1966) );
  AOI22_X1 U1836 ( .A1(n1949), .A2(b[11]), .B1(n1785), .B2(b[10]), .ZN(n1967)
         );
  XNOR2_X1 U1837 ( .A(n1968), .B(n1771), .ZN(n834) );
  OAI221_X1 U1838 ( .B1(n1858), .B2(n1947), .C1(n1853), .C2(n1783), .A(n1969), 
        .ZN(n1968) );
  AOI22_X1 U1839 ( .A1(n1490), .A2(b[12]), .B1(n1471), .B2(b[11]), .ZN(n1969)
         );
  XNOR2_X1 U1840 ( .A(n1970), .B(n1771), .ZN(n833) );
  OAI221_X1 U1841 ( .B1(n1856), .B2(n1947), .C1(n1851), .C2(n1784), .A(n1971), 
        .ZN(n1970) );
  AOI22_X1 U1842 ( .A1(n1490), .A2(b[13]), .B1(n1471), .B2(b[12]), .ZN(n1971)
         );
  XNOR2_X1 U1843 ( .A(n1972), .B(n1770), .ZN(n832) );
  OAI221_X1 U1844 ( .B1(n1854), .B2(n1947), .C1(n1849), .C2(n1783), .A(n1973), 
        .ZN(n1972) );
  AOI22_X1 U1845 ( .A1(n1490), .A2(b[14]), .B1(n1471), .B2(b[13]), .ZN(n1973)
         );
  XNOR2_X1 U1846 ( .A(n1974), .B(n1770), .ZN(n831) );
  OAI221_X1 U1847 ( .B1(n1852), .B2(n1947), .C1(n1632), .C2(n1784), .A(n1975), 
        .ZN(n1974) );
  AOI22_X1 U1848 ( .A1(n1490), .A2(b[15]), .B1(n1471), .B2(b[14]), .ZN(n1975)
         );
  XNOR2_X1 U1849 ( .A(n1976), .B(n1770), .ZN(n830) );
  OAI221_X1 U1850 ( .B1(n1850), .B2(n1947), .C1(n1846), .C2(n1783), .A(n1977), 
        .ZN(n1976) );
  AOI22_X1 U1851 ( .A1(n1490), .A2(b[16]), .B1(n1471), .B2(b[15]), .ZN(n1977)
         );
  XNOR2_X1 U1852 ( .A(n1978), .B(n1770), .ZN(n829) );
  OAI221_X1 U1853 ( .B1(n1848), .B2(n1947), .C1(n1634), .C2(n1783), .A(n1979), 
        .ZN(n1978) );
  AOI22_X1 U1854 ( .A1(n1490), .A2(b[17]), .B1(n1471), .B2(b[16]), .ZN(n1979)
         );
  XNOR2_X1 U1855 ( .A(n1980), .B(n1770), .ZN(n828) );
  OAI221_X1 U1856 ( .B1(n1847), .B2(n1947), .C1(n1843), .C2(n1784), .A(n1981), 
        .ZN(n1980) );
  AOI22_X1 U1857 ( .A1(n1490), .A2(b[18]), .B1(n1471), .B2(b[17]), .ZN(n1981)
         );
  XNOR2_X1 U1858 ( .A(n1982), .B(n1770), .ZN(n827) );
  OAI221_X1 U1859 ( .B1(n1845), .B2(n1947), .C1(n1630), .C2(n1783), .A(n1983), 
        .ZN(n1982) );
  AOI22_X1 U1860 ( .A1(n1490), .A2(b[19]), .B1(n1471), .B2(b[18]), .ZN(n1983)
         );
  XNOR2_X1 U1861 ( .A(n1984), .B(n1770), .ZN(n826) );
  AOI22_X1 U1862 ( .A1(n1490), .A2(b[20]), .B1(n1471), .B2(b[19]), .ZN(n1985)
         );
  XNOR2_X1 U1863 ( .A(n1986), .B(n1770), .ZN(n825) );
  OAI221_X1 U1864 ( .B1(n1842), .B2(n1947), .C1(n1628), .C2(n1783), .A(n1987), 
        .ZN(n1986) );
  AOI22_X1 U1865 ( .A1(n1490), .A2(b[21]), .B1(n1471), .B2(b[20]), .ZN(n1987)
         );
  XNOR2_X1 U1866 ( .A(n1988), .B(n1770), .ZN(n824) );
  AOI22_X1 U1867 ( .A1(n1490), .A2(b[22]), .B1(n1471), .B2(b[21]), .ZN(n1989)
         );
  XNOR2_X1 U1868 ( .A(n1990), .B(n1770), .ZN(n823) );
  OAI21_X1 U1869 ( .B1(n1835), .B2(n1783), .A(n1991), .ZN(n1990) );
  OAI22_X1 U1870 ( .A1(n1824), .A2(n1992), .B1(b[21]), .B2(n1992), .ZN(n1991)
         );
  AOI22_X1 U1871 ( .A1(n1622), .A2(n1588), .B1(n1838), .B2(n1588), .ZN(n1992)
         );
  XNOR2_X1 U1872 ( .A(n1994), .B(n1770), .ZN(n822) );
  OAI21_X1 U1873 ( .B1(n1836), .B2(n1784), .A(n1995), .ZN(n1994) );
  OAI22_X1 U1874 ( .A1(n1824), .A2(n1471), .B1(b[22]), .B2(n1471), .ZN(n1995)
         );
  XNOR2_X1 U1875 ( .A(n1997), .B(n1770), .ZN(n821) );
  OAI21_X1 U1876 ( .B1(n1888), .B2(n1783), .A(n1947), .ZN(n1997) );
  XNOR2_X1 U1877 ( .A(a[6]), .B(a[7]), .ZN(n1996) );
  NAND2_X1 U1878 ( .A1(n1479), .A2(n1993), .ZN(n1944) );
  XNOR2_X1 U1879 ( .A(n1998), .B(n1768), .ZN(n819) );
  OAI22_X1 U1880 ( .A1(n1774), .A2(n1819), .B1(n1775), .B2(n1786), .ZN(n1998)
         );
  XNOR2_X1 U1881 ( .A(n2000), .B(n1769), .ZN(n818) );
  OAI222_X1 U1882 ( .A1(n1775), .A2(n1623), .B1(n1876), .B2(n1819), .C1(n1875), 
        .C2(n1788), .ZN(n2000) );
  XNOR2_X1 U1883 ( .A(n2001), .B(n1769), .ZN(n817) );
  OAI221_X1 U1884 ( .B1(n1774), .B2(n2002), .C1(n1873), .C2(n1787), .A(n2003), 
        .ZN(n2001) );
  AOI22_X1 U1885 ( .A1(n2004), .A2(n1649), .B1(n1789), .B2(n1602), .ZN(n2003)
         );
  XNOR2_X1 U1886 ( .A(n2005), .B(n1769), .ZN(n816) );
  OAI221_X1 U1887 ( .B1(n1876), .B2(n2002), .C1(n1871), .C2(n1787), .A(n2006), 
        .ZN(n2005) );
  AOI22_X1 U1888 ( .A1(n2004), .A2(b[3]), .B1(n1789), .B2(n1649), .ZN(n2006)
         );
  XNOR2_X1 U1889 ( .A(n2007), .B(n1769), .ZN(n815) );
  OAI221_X1 U1890 ( .B1(n1874), .B2(n2002), .C1(n1869), .C2(n1787), .A(n2008), 
        .ZN(n2007) );
  AOI22_X1 U1891 ( .A1(n2004), .A2(b[4]), .B1(n1789), .B2(b[3]), .ZN(n2008) );
  XNOR2_X1 U1892 ( .A(n2009), .B(n1769), .ZN(n814) );
  OAI221_X1 U1893 ( .B1(n1872), .B2(n2002), .C1(n1867), .C2(n1787), .A(n2010), 
        .ZN(n2009) );
  AOI22_X1 U1894 ( .A1(n2004), .A2(b[5]), .B1(n1789), .B2(b[4]), .ZN(n2010) );
  XNOR2_X1 U1895 ( .A(n2011), .B(n1769), .ZN(n813) );
  OAI221_X1 U1896 ( .B1(n1870), .B2(n2002), .C1(n1865), .C2(n1787), .A(n2012), 
        .ZN(n2011) );
  AOI22_X1 U1897 ( .A1(n2004), .A2(b[6]), .B1(n1789), .B2(b[5]), .ZN(n2012) );
  XNOR2_X1 U1898 ( .A(n2013), .B(n1769), .ZN(n812) );
  OAI221_X1 U1899 ( .B1(n1868), .B2(n2002), .C1(n1863), .C2(n1787), .A(n2014), 
        .ZN(n2013) );
  AOI22_X1 U1900 ( .A1(n2004), .A2(b[7]), .B1(n1789), .B2(b[6]), .ZN(n2014) );
  XNOR2_X1 U1901 ( .A(n2015), .B(n1769), .ZN(n811) );
  OAI221_X1 U1902 ( .B1(n1866), .B2(n2002), .C1(n1861), .C2(n1787), .A(n2016), 
        .ZN(n2015) );
  AOI22_X1 U1903 ( .A1(n2004), .A2(b[8]), .B1(n1789), .B2(b[7]), .ZN(n2016) );
  XNOR2_X1 U1904 ( .A(n2017), .B(n1769), .ZN(n810) );
  OAI221_X1 U1905 ( .B1(n1864), .B2(n2002), .C1(n1859), .C2(n1787), .A(n2018), 
        .ZN(n2017) );
  AOI22_X1 U1906 ( .A1(n2004), .A2(b[9]), .B1(n1789), .B2(b[8]), .ZN(n2018) );
  XNOR2_X1 U1907 ( .A(n2019), .B(n1769), .ZN(n809) );
  OAI221_X1 U1908 ( .B1(n1862), .B2(n2002), .C1(n1857), .C2(n1787), .A(n2020), 
        .ZN(n2019) );
  AOI22_X1 U1909 ( .A1(n2004), .A2(b[10]), .B1(n1789), .B2(b[9]), .ZN(n2020)
         );
  XNOR2_X1 U1910 ( .A(n2021), .B(n1769), .ZN(n808) );
  OAI221_X1 U1911 ( .B1(n1860), .B2(n2002), .C1(n1855), .C2(n1787), .A(n2022), 
        .ZN(n2021) );
  AOI22_X1 U1912 ( .A1(n2004), .A2(b[11]), .B1(n1789), .B2(b[10]), .ZN(n2022)
         );
  XNOR2_X1 U1913 ( .A(n2023), .B(n1769), .ZN(n807) );
  OAI221_X1 U1914 ( .B1(n1858), .B2(n2002), .C1(n1853), .C2(n1786), .A(n2024), 
        .ZN(n2023) );
  AOI22_X1 U1915 ( .A1(n2004), .A2(b[12]), .B1(n1789), .B2(b[11]), .ZN(n2024)
         );
  XNOR2_X1 U1916 ( .A(n2025), .B(n1769), .ZN(n806) );
  OAI221_X1 U1917 ( .B1(n1856), .B2(n2002), .C1(n1851), .C2(n1786), .A(n2026), 
        .ZN(n2025) );
  AOI22_X1 U1918 ( .A1(n2004), .A2(b[13]), .B1(n1789), .B2(b[12]), .ZN(n2026)
         );
  XNOR2_X1 U1919 ( .A(n2027), .B(n1768), .ZN(n805) );
  OAI221_X1 U1920 ( .B1(n1854), .B2(n2002), .C1(n1849), .C2(n1786), .A(n2028), 
        .ZN(n2027) );
  AOI22_X1 U1921 ( .A1(n2004), .A2(b[14]), .B1(n1789), .B2(b[13]), .ZN(n2028)
         );
  XNOR2_X1 U1922 ( .A(n2029), .B(n1768), .ZN(n804) );
  OAI221_X1 U1923 ( .B1(n1852), .B2(n2002), .C1(n1632), .C2(n1786), .A(n2030), 
        .ZN(n2029) );
  AOI22_X1 U1924 ( .A1(n2004), .A2(b[15]), .B1(n1789), .B2(b[14]), .ZN(n2030)
         );
  XNOR2_X1 U1925 ( .A(n2031), .B(n1768), .ZN(n803) );
  OAI221_X1 U1926 ( .B1(n1850), .B2(n2002), .C1(n1846), .C2(n1786), .A(n2032), 
        .ZN(n2031) );
  AOI22_X1 U1927 ( .A1(n2004), .A2(b[16]), .B1(n1789), .B2(b[15]), .ZN(n2032)
         );
  XNOR2_X1 U1928 ( .A(n2033), .B(n1768), .ZN(n802) );
  AOI22_X1 U1929 ( .A1(n2004), .A2(b[17]), .B1(n1789), .B2(b[16]), .ZN(n2034)
         );
  XNOR2_X1 U1930 ( .A(n2035), .B(n1768), .ZN(n801) );
  OAI221_X1 U1931 ( .B1(n1847), .B2(n2002), .C1(n1843), .C2(n1786), .A(n2036), 
        .ZN(n2035) );
  AOI22_X1 U1932 ( .A1(n2004), .A2(b[18]), .B1(n1789), .B2(b[17]), .ZN(n2036)
         );
  XNOR2_X1 U1933 ( .A(n2037), .B(n1768), .ZN(n800) );
  OAI221_X1 U1934 ( .B1(n1845), .B2(n2002), .C1(n1486), .C2(n1786), .A(n2038), 
        .ZN(n2037) );
  AOI22_X1 U1935 ( .A1(n2004), .A2(b[19]), .B1(n1789), .B2(b[18]), .ZN(n2038)
         );
  XNOR2_X1 U1936 ( .A(n2039), .B(n1768), .ZN(n799) );
  OAI221_X1 U1937 ( .B1(n1844), .B2(n2002), .C1(n1840), .C2(n1786), .A(n2040), 
        .ZN(n2039) );
  AOI22_X1 U1938 ( .A1(n2004), .A2(b[20]), .B1(n1789), .B2(b[19]), .ZN(n2040)
         );
  XNOR2_X1 U1939 ( .A(n2041), .B(n1768), .ZN(n798) );
  OAI221_X1 U1940 ( .B1(n1842), .B2(n2002), .C1(n1628), .C2(n1786), .A(n2042), 
        .ZN(n2041) );
  AOI22_X1 U1941 ( .A1(n2004), .A2(b[21]), .B1(n1789), .B2(b[20]), .ZN(n2042)
         );
  XNOR2_X1 U1942 ( .A(n2043), .B(n1768), .ZN(n797) );
  AOI22_X1 U1943 ( .A1(n2004), .A2(b[22]), .B1(n1789), .B2(b[21]), .ZN(n2044)
         );
  XNOR2_X1 U1944 ( .A(n2045), .B(n1768), .ZN(n796) );
  OAI21_X1 U1945 ( .B1(n1835), .B2(n1787), .A(n2046), .ZN(n2045) );
  OAI22_X1 U1946 ( .A1(n1818), .A2(n2047), .B1(b[21]), .B2(n2047), .ZN(n2046)
         );
  AOI22_X1 U1947 ( .A1(n1623), .A2(n1819), .B1(n1838), .B2(n1819), .ZN(n2047)
         );
  XNOR2_X1 U1948 ( .A(n2050), .B(n1768), .ZN(n795) );
  OAI21_X1 U1949 ( .B1(n1836), .B2(n1788), .A(n2051), .ZN(n2050) );
  OAI22_X1 U1950 ( .A1(n1818), .A2(n1789), .B1(b[22]), .B2(n1789), .ZN(n2051)
         );
  XNOR2_X1 U1951 ( .A(n2053), .B(n1768), .ZN(n794) );
  OAI21_X1 U1952 ( .B1(n1888), .B2(n1787), .A(n2002), .ZN(n2053) );
  XNOR2_X1 U1953 ( .A(a[10]), .B(a[9]), .ZN(n2052) );
  NAND2_X1 U1954 ( .A1(n1821), .A2(n2048), .ZN(n1999) );
  XNOR2_X1 U1955 ( .A(a[10]), .B(n1768), .ZN(n2048) );
  XNOR2_X1 U1956 ( .A(n2054), .B(n1766), .ZN(n792) );
  OAI22_X1 U1957 ( .A1(n1774), .A2(n1813), .B1(n1775), .B2(n1790), .ZN(n2054)
         );
  XNOR2_X1 U1958 ( .A(n2055), .B(n1767), .ZN(n791) );
  OAI222_X1 U1959 ( .A1(n1775), .A2(n1815), .B1(n1876), .B2(n1813), .C1(n1875), 
        .C2(n1790), .ZN(n2055) );
  XNOR2_X1 U1960 ( .A(n2056), .B(n1767), .ZN(n790) );
  OAI221_X1 U1961 ( .B1(n1774), .B2(n2057), .C1(n1873), .C2(n1790), .A(n2058), 
        .ZN(n2056) );
  AOI22_X1 U1962 ( .A1(n2059), .A2(n1649), .B1(n2060), .B2(n1602), .ZN(n2058)
         );
  XNOR2_X1 U1963 ( .A(n2061), .B(n1767), .ZN(n789) );
  OAI221_X1 U1964 ( .B1(n1876), .B2(n2057), .C1(n1871), .C2(n1790), .A(n2062), 
        .ZN(n2061) );
  AOI22_X1 U1965 ( .A1(n2059), .A2(b[3]), .B1(n2060), .B2(n1649), .ZN(n2062)
         );
  XNOR2_X1 U1966 ( .A(n2063), .B(n1767), .ZN(n788) );
  OAI221_X1 U1967 ( .B1(n1874), .B2(n2057), .C1(n1869), .C2(n1790), .A(n2064), 
        .ZN(n2063) );
  AOI22_X1 U1968 ( .A1(n2059), .A2(b[4]), .B1(n2060), .B2(b[3]), .ZN(n2064) );
  XNOR2_X1 U1969 ( .A(n2065), .B(n1767), .ZN(n787) );
  OAI221_X1 U1970 ( .B1(n1872), .B2(n2057), .C1(n1867), .C2(n1790), .A(n2066), 
        .ZN(n2065) );
  AOI22_X1 U1971 ( .A1(n2059), .A2(b[5]), .B1(n2060), .B2(b[4]), .ZN(n2066) );
  XNOR2_X1 U1972 ( .A(n2067), .B(n1767), .ZN(n786) );
  OAI221_X1 U1973 ( .B1(n1870), .B2(n2057), .C1(n1865), .C2(n1790), .A(n2068), 
        .ZN(n2067) );
  AOI22_X1 U1974 ( .A1(n2059), .A2(b[6]), .B1(n2060), .B2(b[5]), .ZN(n2068) );
  XNOR2_X1 U1975 ( .A(n2069), .B(n1767), .ZN(n785) );
  OAI221_X1 U1976 ( .B1(n1868), .B2(n2057), .C1(n1863), .C2(n1790), .A(n2070), 
        .ZN(n2069) );
  AOI22_X1 U1977 ( .A1(n2059), .A2(b[7]), .B1(n2060), .B2(b[6]), .ZN(n2070) );
  XNOR2_X1 U1978 ( .A(n2071), .B(n1767), .ZN(n784) );
  OAI221_X1 U1979 ( .B1(n1866), .B2(n2057), .C1(n1861), .C2(n1790), .A(n2072), 
        .ZN(n2071) );
  AOI22_X1 U1980 ( .A1(n2059), .A2(b[8]), .B1(n2060), .B2(b[7]), .ZN(n2072) );
  XNOR2_X1 U1981 ( .A(n2073), .B(n1767), .ZN(n783) );
  OAI221_X1 U1982 ( .B1(n1864), .B2(n2057), .C1(n1859), .C2(n1790), .A(n2074), 
        .ZN(n2073) );
  AOI22_X1 U1983 ( .A1(n2059), .A2(b[9]), .B1(n2060), .B2(b[8]), .ZN(n2074) );
  XNOR2_X1 U1984 ( .A(n2075), .B(n1767), .ZN(n782) );
  OAI221_X1 U1985 ( .B1(n1862), .B2(n2057), .C1(n1857), .C2(n1790), .A(n2076), 
        .ZN(n2075) );
  AOI22_X1 U1986 ( .A1(n2059), .A2(b[10]), .B1(n2060), .B2(b[9]), .ZN(n2076)
         );
  XNOR2_X1 U1987 ( .A(n2077), .B(n1767), .ZN(n781) );
  OAI221_X1 U1988 ( .B1(n1860), .B2(n2057), .C1(n1855), .C2(n1790), .A(n2078), 
        .ZN(n2077) );
  AOI22_X1 U1989 ( .A1(n2059), .A2(b[11]), .B1(n2060), .B2(b[10]), .ZN(n2078)
         );
  XNOR2_X1 U1990 ( .A(n2079), .B(n1767), .ZN(n780) );
  OAI221_X1 U1991 ( .B1(n1858), .B2(n2057), .C1(n1853), .C2(n1790), .A(n2080), 
        .ZN(n2079) );
  AOI22_X1 U1992 ( .A1(n2059), .A2(b[12]), .B1(n2060), .B2(b[11]), .ZN(n2080)
         );
  XNOR2_X1 U1993 ( .A(n2081), .B(n1766), .ZN(n779) );
  OAI221_X1 U1994 ( .B1(n1856), .B2(n2057), .C1(n1851), .C2(n1790), .A(n2082), 
        .ZN(n2081) );
  AOI22_X1 U1995 ( .A1(n2059), .A2(b[13]), .B1(n2060), .B2(b[12]), .ZN(n2082)
         );
  XNOR2_X1 U1996 ( .A(n2083), .B(n1766), .ZN(n778) );
  OAI221_X1 U1997 ( .B1(n1854), .B2(n2057), .C1(n1849), .C2(n1790), .A(n2084), 
        .ZN(n2083) );
  AOI22_X1 U1998 ( .A1(n2059), .A2(b[14]), .B1(n2060), .B2(b[13]), .ZN(n2084)
         );
  XNOR2_X1 U1999 ( .A(n2085), .B(n1766), .ZN(n777) );
  OAI221_X1 U2000 ( .B1(n1852), .B2(n2057), .C1(n1632), .C2(n1790), .A(n2086), 
        .ZN(n2085) );
  AOI22_X1 U2001 ( .A1(n2059), .A2(b[15]), .B1(n2060), .B2(b[14]), .ZN(n2086)
         );
  XNOR2_X1 U2002 ( .A(n2087), .B(n1766), .ZN(n776) );
  OAI221_X1 U2003 ( .B1(n1850), .B2(n2057), .C1(n1846), .C2(n1790), .A(n2088), 
        .ZN(n2087) );
  AOI22_X1 U2004 ( .A1(n2059), .A2(b[16]), .B1(n2060), .B2(b[15]), .ZN(n2088)
         );
  XNOR2_X1 U2005 ( .A(n2089), .B(n1766), .ZN(n775) );
  AOI22_X1 U2006 ( .A1(n2059), .A2(b[17]), .B1(n2060), .B2(b[16]), .ZN(n2090)
         );
  XNOR2_X1 U2007 ( .A(n2091), .B(n1766), .ZN(n774) );
  OAI221_X1 U2008 ( .B1(n1847), .B2(n2057), .C1(n1843), .C2(n1790), .A(n2092), 
        .ZN(n2091) );
  AOI22_X1 U2009 ( .A1(n2059), .A2(b[18]), .B1(n2060), .B2(b[17]), .ZN(n2092)
         );
  XNOR2_X1 U2010 ( .A(n2093), .B(n1766), .ZN(n773) );
  OAI221_X1 U2011 ( .B1(n1845), .B2(n2057), .C1(n1493), .C2(n1790), .A(n2094), 
        .ZN(n2093) );
  AOI22_X1 U2012 ( .A1(n2059), .A2(b[19]), .B1(n2060), .B2(b[18]), .ZN(n2094)
         );
  XNOR2_X1 U2013 ( .A(n2095), .B(n1766), .ZN(n772) );
  OAI221_X1 U2014 ( .B1(n1844), .B2(n2057), .C1(n1840), .C2(n1790), .A(n2096), 
        .ZN(n2095) );
  AOI22_X1 U2015 ( .A1(n2059), .A2(b[20]), .B1(n2060), .B2(b[19]), .ZN(n2096)
         );
  XNOR2_X1 U2016 ( .A(n2097), .B(n1766), .ZN(n771) );
  OAI221_X1 U2017 ( .B1(n1842), .B2(n2057), .C1(n1494), .C2(n1790), .A(n2098), 
        .ZN(n2097) );
  AOI22_X1 U2018 ( .A1(n2059), .A2(b[21]), .B1(n2060), .B2(b[20]), .ZN(n2098)
         );
  XNOR2_X1 U2019 ( .A(a[14]), .B(n2099), .ZN(n770) );
  AOI221_X1 U2020 ( .B1(n2059), .B2(b[22]), .C1(n1472), .C2(n1497), .A(n2100), 
        .ZN(n2099) );
  OAI22_X1 U2021 ( .A1(n1841), .A2(n2057), .B1(n1839), .B2(n1815), .ZN(n2100)
         );
  XNOR2_X1 U2022 ( .A(n2101), .B(n1766), .ZN(n769) );
  OAI21_X1 U2023 ( .B1(n1835), .B2(n1790), .A(n2102), .ZN(n2101) );
  OAI22_X1 U2024 ( .A1(n1812), .A2(n2103), .B1(b[21]), .B2(n2103), .ZN(n2102)
         );
  AOI22_X1 U2025 ( .A1(n1815), .A2(n1813), .B1(n1838), .B2(n1813), .ZN(n2103)
         );
  XNOR2_X1 U2026 ( .A(n2106), .B(n1766), .ZN(n768) );
  OAI21_X1 U2027 ( .B1(n1836), .B2(n1790), .A(n2107), .ZN(n2106) );
  OAI22_X1 U2028 ( .A1(n1812), .A2(n2060), .B1(b[22]), .B2(n2060), .ZN(n2107)
         );
  XNOR2_X1 U2029 ( .A(n2109), .B(n1766), .ZN(n767) );
  OAI21_X1 U2030 ( .B1(n1888), .B2(n1790), .A(n2057), .ZN(n2109) );
  XNOR2_X1 U2031 ( .A(a[12]), .B(a[13]), .ZN(n2108) );
  XNOR2_X1 U2032 ( .A(a[13]), .B(n1766), .ZN(n2104) );
  XOR2_X1 U2033 ( .A(a[12]), .B(n1820), .Z(n2105) );
  XNOR2_X1 U2034 ( .A(n2110), .B(n1764), .ZN(n765) );
  OAI22_X1 U2035 ( .A1(n1774), .A2(n1808), .B1(n1775), .B2(n1791), .ZN(n2110)
         );
  XNOR2_X1 U2036 ( .A(n2111), .B(n1765), .ZN(n764) );
  OAI222_X1 U2037 ( .A1(n1775), .A2(n1810), .B1(n1876), .B2(n1808), .C1(n1875), 
        .C2(n1791), .ZN(n2111) );
  XNOR2_X1 U2038 ( .A(n2112), .B(n1765), .ZN(n763) );
  OAI221_X1 U2039 ( .B1(n1774), .B2(n2113), .C1(n1873), .C2(n1791), .A(n2114), 
        .ZN(n2112) );
  AOI22_X1 U2040 ( .A1(n2115), .A2(n1649), .B1(n2116), .B2(n1745), .ZN(n2114)
         );
  XNOR2_X1 U2041 ( .A(n2117), .B(n1765), .ZN(n762) );
  OAI221_X1 U2042 ( .B1(n1876), .B2(n2113), .C1(n1871), .C2(n1791), .A(n2118), 
        .ZN(n2117) );
  AOI22_X1 U2043 ( .A1(n2115), .A2(b[3]), .B1(n2116), .B2(n1649), .ZN(n2118)
         );
  XNOR2_X1 U2044 ( .A(n2119), .B(n1765), .ZN(n761) );
  OAI221_X1 U2045 ( .B1(n1874), .B2(n2113), .C1(n1869), .C2(n1791), .A(n2120), 
        .ZN(n2119) );
  AOI22_X1 U2046 ( .A1(n2115), .A2(b[4]), .B1(n2116), .B2(b[3]), .ZN(n2120) );
  XNOR2_X1 U2047 ( .A(n2121), .B(n1765), .ZN(n760) );
  OAI221_X1 U2048 ( .B1(n1872), .B2(n2113), .C1(n1867), .C2(n1791), .A(n2122), 
        .ZN(n2121) );
  AOI22_X1 U2049 ( .A1(n2115), .A2(b[5]), .B1(n2116), .B2(b[4]), .ZN(n2122) );
  XNOR2_X1 U2050 ( .A(n2123), .B(n1765), .ZN(n759) );
  OAI221_X1 U2051 ( .B1(n1870), .B2(n2113), .C1(n1865), .C2(n1791), .A(n2124), 
        .ZN(n2123) );
  AOI22_X1 U2052 ( .A1(n2115), .A2(b[6]), .B1(n2116), .B2(b[5]), .ZN(n2124) );
  XNOR2_X1 U2053 ( .A(n2125), .B(n1765), .ZN(n758) );
  OAI221_X1 U2054 ( .B1(n1868), .B2(n2113), .C1(n1863), .C2(n1791), .A(n2126), 
        .ZN(n2125) );
  AOI22_X1 U2055 ( .A1(n2115), .A2(b[7]), .B1(n2116), .B2(b[6]), .ZN(n2126) );
  XNOR2_X1 U2056 ( .A(n2127), .B(n1765), .ZN(n757) );
  OAI221_X1 U2057 ( .B1(n1866), .B2(n2113), .C1(n1861), .C2(n1791), .A(n2128), 
        .ZN(n2127) );
  AOI22_X1 U2058 ( .A1(n2115), .A2(b[8]), .B1(n2116), .B2(b[7]), .ZN(n2128) );
  XNOR2_X1 U2059 ( .A(n2129), .B(n1765), .ZN(n756) );
  OAI221_X1 U2060 ( .B1(n1864), .B2(n2113), .C1(n1859), .C2(n1791), .A(n2130), 
        .ZN(n2129) );
  AOI22_X1 U2061 ( .A1(n2115), .A2(b[9]), .B1(n2116), .B2(b[8]), .ZN(n2130) );
  XNOR2_X1 U2062 ( .A(n2131), .B(n1765), .ZN(n755) );
  OAI221_X1 U2063 ( .B1(n1862), .B2(n2113), .C1(n1857), .C2(n1791), .A(n2132), 
        .ZN(n2131) );
  AOI22_X1 U2064 ( .A1(n2115), .A2(b[10]), .B1(n2116), .B2(b[9]), .ZN(n2132)
         );
  XNOR2_X1 U2065 ( .A(n2133), .B(n1765), .ZN(n754) );
  OAI221_X1 U2066 ( .B1(n1860), .B2(n2113), .C1(n1855), .C2(n1791), .A(n2134), 
        .ZN(n2133) );
  AOI22_X1 U2067 ( .A1(n2115), .A2(b[11]), .B1(n2116), .B2(b[10]), .ZN(n2134)
         );
  XNOR2_X1 U2068 ( .A(n2135), .B(n1765), .ZN(n753) );
  OAI221_X1 U2069 ( .B1(n1858), .B2(n2113), .C1(n1853), .C2(n1791), .A(n2136), 
        .ZN(n2135) );
  AOI22_X1 U2070 ( .A1(n2115), .A2(b[12]), .B1(n2116), .B2(b[11]), .ZN(n2136)
         );
  XNOR2_X1 U2071 ( .A(n2137), .B(n1764), .ZN(n752) );
  OAI221_X1 U2072 ( .B1(n1856), .B2(n2113), .C1(n1851), .C2(n1791), .A(n2138), 
        .ZN(n2137) );
  AOI22_X1 U2073 ( .A1(n2115), .A2(b[13]), .B1(n2116), .B2(b[12]), .ZN(n2138)
         );
  XNOR2_X1 U2074 ( .A(n2139), .B(n1764), .ZN(n751) );
  OAI221_X1 U2075 ( .B1(n1854), .B2(n2113), .C1(n1849), .C2(n1791), .A(n2140), 
        .ZN(n2139) );
  AOI22_X1 U2076 ( .A1(n2115), .A2(b[14]), .B1(n2116), .B2(b[13]), .ZN(n2140)
         );
  XNOR2_X1 U2077 ( .A(n2141), .B(n1764), .ZN(n750) );
  OAI221_X1 U2078 ( .B1(n1852), .B2(n2113), .C1(n1632), .C2(n1791), .A(n2142), 
        .ZN(n2141) );
  AOI22_X1 U2079 ( .A1(n2115), .A2(b[15]), .B1(n2116), .B2(b[14]), .ZN(n2142)
         );
  XNOR2_X1 U2080 ( .A(n2143), .B(n1764), .ZN(n749) );
  OAI221_X1 U2081 ( .B1(n1850), .B2(n2113), .C1(n1846), .C2(n1791), .A(n2144), 
        .ZN(n2143) );
  AOI22_X1 U2082 ( .A1(n2115), .A2(b[16]), .B1(n2116), .B2(b[15]), .ZN(n2144)
         );
  XNOR2_X1 U2083 ( .A(n2145), .B(n1764), .ZN(n748) );
  AOI22_X1 U2084 ( .A1(n2115), .A2(b[17]), .B1(n2116), .B2(b[16]), .ZN(n2146)
         );
  XNOR2_X1 U2085 ( .A(n2147), .B(n1764), .ZN(n747) );
  OAI221_X1 U2086 ( .B1(n1847), .B2(n2113), .C1(n1843), .C2(n1791), .A(n2148), 
        .ZN(n2147) );
  AOI22_X1 U2087 ( .A1(n2115), .A2(b[18]), .B1(n2116), .B2(b[17]), .ZN(n2148)
         );
  XNOR2_X1 U2088 ( .A(n2149), .B(n1764), .ZN(n746) );
  OAI221_X1 U2089 ( .B1(n1845), .B2(n2113), .C1(n1493), .C2(n1791), .A(n2150), 
        .ZN(n2149) );
  AOI22_X1 U2090 ( .A1(n2115), .A2(b[19]), .B1(n2116), .B2(b[18]), .ZN(n2150)
         );
  XNOR2_X1 U2091 ( .A(n2151), .B(n1764), .ZN(n745) );
  OAI221_X1 U2092 ( .B1(n1844), .B2(n2113), .C1(n1840), .C2(n1791), .A(n2152), 
        .ZN(n2151) );
  AOI22_X1 U2093 ( .A1(n2115), .A2(b[20]), .B1(n2116), .B2(b[19]), .ZN(n2152)
         );
  XNOR2_X1 U2094 ( .A(n2153), .B(n1764), .ZN(n744) );
  OAI221_X1 U2095 ( .B1(n1842), .B2(n2113), .C1(n1494), .C2(n1791), .A(n2154), 
        .ZN(n2153) );
  AOI22_X1 U2096 ( .A1(n2115), .A2(b[21]), .B1(n2116), .B2(b[20]), .ZN(n2154)
         );
  XNOR2_X1 U2097 ( .A(a[17]), .B(n2155), .ZN(n743) );
  AOI221_X1 U2098 ( .B1(n2115), .B2(b[22]), .C1(n1621), .C2(n1497), .A(n2156), 
        .ZN(n2155) );
  OAI22_X1 U2099 ( .A1(n1841), .A2(n2113), .B1(n1839), .B2(n1810), .ZN(n2156)
         );
  XNOR2_X1 U2100 ( .A(n2157), .B(n1764), .ZN(n742) );
  OAI21_X1 U2101 ( .B1(n1835), .B2(n1791), .A(n2158), .ZN(n2157) );
  OAI22_X1 U2102 ( .A1(n1807), .A2(n2159), .B1(b[21]), .B2(n2159), .ZN(n2158)
         );
  AOI22_X1 U2103 ( .A1(n1810), .A2(n1808), .B1(n1838), .B2(n1808), .ZN(n2159)
         );
  XNOR2_X1 U2104 ( .A(n2162), .B(n1764), .ZN(n741) );
  OAI21_X1 U2105 ( .B1(n1836), .B2(n1791), .A(n2163), .ZN(n2162) );
  OAI22_X1 U2106 ( .A1(n1807), .A2(n2116), .B1(b[22]), .B2(n2116), .ZN(n2163)
         );
  XNOR2_X1 U2107 ( .A(n2165), .B(n1764), .ZN(n740) );
  OAI21_X1 U2108 ( .B1(n1888), .B2(n1791), .A(n2113), .ZN(n2165) );
  XNOR2_X1 U2109 ( .A(a[15]), .B(a[16]), .ZN(n2164) );
  XNOR2_X1 U2110 ( .A(a[16]), .B(n1764), .ZN(n2160) );
  XOR2_X1 U2111 ( .A(a[15]), .B(n1767), .Z(n2161) );
  XNOR2_X1 U2112 ( .A(n2166), .B(n1762), .ZN(n738) );
  OAI22_X1 U2113 ( .A1(n1774), .A2(n1803), .B1(n1775), .B2(n1792), .ZN(n2166)
         );
  XNOR2_X1 U2114 ( .A(n2167), .B(n1763), .ZN(n737) );
  OAI222_X1 U2115 ( .A1(n1775), .A2(n1805), .B1(n1876), .B2(n1803), .C1(n1875), 
        .C2(n1792), .ZN(n2167) );
  XNOR2_X1 U2116 ( .A(n2168), .B(n1763), .ZN(n736) );
  OAI221_X1 U2117 ( .B1(n1774), .B2(n2169), .C1(n1873), .C2(n1792), .A(n2170), 
        .ZN(n2168) );
  AOI22_X1 U2118 ( .A1(n2171), .A2(n1649), .B1(n2172), .B2(n1745), .ZN(n2170)
         );
  XNOR2_X1 U2119 ( .A(n2173), .B(n1763), .ZN(n735) );
  OAI221_X1 U2120 ( .B1(n1876), .B2(n2169), .C1(n1871), .C2(n1792), .A(n2174), 
        .ZN(n2173) );
  AOI22_X1 U2121 ( .A1(n2171), .A2(b[3]), .B1(n2172), .B2(n1649), .ZN(n2174)
         );
  XNOR2_X1 U2122 ( .A(n2175), .B(n1763), .ZN(n734) );
  OAI221_X1 U2123 ( .B1(n1874), .B2(n2169), .C1(n1869), .C2(n1792), .A(n2176), 
        .ZN(n2175) );
  AOI22_X1 U2124 ( .A1(n2171), .A2(b[4]), .B1(n2172), .B2(b[3]), .ZN(n2176) );
  XNOR2_X1 U2125 ( .A(n2177), .B(n1763), .ZN(n733) );
  OAI221_X1 U2126 ( .B1(n1872), .B2(n2169), .C1(n1867), .C2(n1792), .A(n2178), 
        .ZN(n2177) );
  AOI22_X1 U2127 ( .A1(n2171), .A2(b[5]), .B1(n2172), .B2(b[4]), .ZN(n2178) );
  XNOR2_X1 U2128 ( .A(n2179), .B(n1763), .ZN(n732) );
  OAI221_X1 U2129 ( .B1(n1870), .B2(n2169), .C1(n1865), .C2(n1792), .A(n2180), 
        .ZN(n2179) );
  AOI22_X1 U2130 ( .A1(n2171), .A2(b[6]), .B1(n2172), .B2(b[5]), .ZN(n2180) );
  XNOR2_X1 U2131 ( .A(n2181), .B(n1763), .ZN(n731) );
  OAI221_X1 U2132 ( .B1(n1868), .B2(n2169), .C1(n1863), .C2(n1792), .A(n2182), 
        .ZN(n2181) );
  AOI22_X1 U2133 ( .A1(n2171), .A2(b[7]), .B1(n2172), .B2(b[6]), .ZN(n2182) );
  XNOR2_X1 U2134 ( .A(n2183), .B(n1763), .ZN(n730) );
  OAI221_X1 U2135 ( .B1(n1866), .B2(n2169), .C1(n1861), .C2(n1792), .A(n2184), 
        .ZN(n2183) );
  AOI22_X1 U2136 ( .A1(n2171), .A2(b[8]), .B1(n2172), .B2(b[7]), .ZN(n2184) );
  XNOR2_X1 U2137 ( .A(n2185), .B(n1763), .ZN(n729) );
  OAI221_X1 U2138 ( .B1(n1864), .B2(n2169), .C1(n1859), .C2(n1792), .A(n2186), 
        .ZN(n2185) );
  AOI22_X1 U2139 ( .A1(n2171), .A2(b[9]), .B1(n2172), .B2(b[8]), .ZN(n2186) );
  XNOR2_X1 U2140 ( .A(n2187), .B(n1763), .ZN(n728) );
  OAI221_X1 U2141 ( .B1(n1862), .B2(n2169), .C1(n1857), .C2(n1792), .A(n2188), 
        .ZN(n2187) );
  AOI22_X1 U2142 ( .A1(n2171), .A2(b[10]), .B1(n2172), .B2(b[9]), .ZN(n2188)
         );
  XNOR2_X1 U2143 ( .A(n2189), .B(n1763), .ZN(n727) );
  OAI221_X1 U2144 ( .B1(n1860), .B2(n2169), .C1(n1855), .C2(n1792), .A(n2190), 
        .ZN(n2189) );
  AOI22_X1 U2145 ( .A1(n2171), .A2(b[11]), .B1(n2172), .B2(b[10]), .ZN(n2190)
         );
  XNOR2_X1 U2146 ( .A(n2191), .B(n1763), .ZN(n726) );
  OAI221_X1 U2147 ( .B1(n1858), .B2(n2169), .C1(n1853), .C2(n1792), .A(n2192), 
        .ZN(n2191) );
  AOI22_X1 U2148 ( .A1(n2171), .A2(b[12]), .B1(n2172), .B2(b[11]), .ZN(n2192)
         );
  XNOR2_X1 U2149 ( .A(n2193), .B(n1762), .ZN(n725) );
  OAI221_X1 U2150 ( .B1(n1856), .B2(n2169), .C1(n1851), .C2(n1792), .A(n2194), 
        .ZN(n2193) );
  AOI22_X1 U2151 ( .A1(n2171), .A2(b[13]), .B1(n2172), .B2(b[12]), .ZN(n2194)
         );
  XNOR2_X1 U2152 ( .A(n2195), .B(n1762), .ZN(n724) );
  OAI221_X1 U2153 ( .B1(n1854), .B2(n2169), .C1(n1849), .C2(n1792), .A(n2196), 
        .ZN(n2195) );
  AOI22_X1 U2154 ( .A1(n2171), .A2(b[14]), .B1(n2172), .B2(b[13]), .ZN(n2196)
         );
  XNOR2_X1 U2155 ( .A(n2197), .B(n1762), .ZN(n723) );
  OAI221_X1 U2156 ( .B1(n1852), .B2(n2169), .C1(n1632), .C2(n1792), .A(n2198), 
        .ZN(n2197) );
  AOI22_X1 U2157 ( .A1(n2171), .A2(b[15]), .B1(n2172), .B2(b[14]), .ZN(n2198)
         );
  XNOR2_X1 U2158 ( .A(n2199), .B(n1762), .ZN(n722) );
  OAI221_X1 U2159 ( .B1(n1850), .B2(n2169), .C1(n1846), .C2(n1792), .A(n2200), 
        .ZN(n2199) );
  AOI22_X1 U2160 ( .A1(n2171), .A2(b[16]), .B1(n2172), .B2(b[15]), .ZN(n2200)
         );
  XNOR2_X1 U2161 ( .A(n2201), .B(n1762), .ZN(n721) );
  AOI22_X1 U2162 ( .A1(n2171), .A2(b[17]), .B1(n2172), .B2(b[16]), .ZN(n2202)
         );
  XNOR2_X1 U2163 ( .A(n2203), .B(n1762), .ZN(n720) );
  OAI221_X1 U2164 ( .B1(n1847), .B2(n2169), .C1(n1843), .C2(n1792), .A(n2204), 
        .ZN(n2203) );
  AOI22_X1 U2165 ( .A1(n2171), .A2(b[18]), .B1(n2172), .B2(b[17]), .ZN(n2204)
         );
  XNOR2_X1 U2166 ( .A(n2205), .B(n1762), .ZN(n719) );
  OAI221_X1 U2167 ( .B1(n1845), .B2(n2169), .C1(n1493), .C2(n1792), .A(n2206), 
        .ZN(n2205) );
  AOI22_X1 U2168 ( .A1(n2171), .A2(b[19]), .B1(n2172), .B2(b[18]), .ZN(n2206)
         );
  XNOR2_X1 U2169 ( .A(n2207), .B(n1762), .ZN(n718) );
  OAI221_X1 U2170 ( .B1(n1844), .B2(n2169), .C1(n1840), .C2(n1792), .A(n2208), 
        .ZN(n2207) );
  AOI22_X1 U2171 ( .A1(n2171), .A2(b[20]), .B1(n2172), .B2(b[19]), .ZN(n2208)
         );
  XNOR2_X1 U2172 ( .A(n2209), .B(n1762), .ZN(n717) );
  OAI221_X1 U2173 ( .B1(n1842), .B2(n2169), .C1(n1494), .C2(n1792), .A(n2210), 
        .ZN(n2209) );
  AOI22_X1 U2174 ( .A1(n2171), .A2(b[21]), .B1(n2172), .B2(b[20]), .ZN(n2210)
         );
  XNOR2_X1 U2175 ( .A(a[20]), .B(n2211), .ZN(n716) );
  OAI22_X1 U2176 ( .A1(n1841), .A2(n2169), .B1(n1839), .B2(n1805), .ZN(n2212)
         );
  XNOR2_X1 U2177 ( .A(n2213), .B(n1762), .ZN(n715) );
  OAI21_X1 U2178 ( .B1(n1835), .B2(n1792), .A(n2214), .ZN(n2213) );
  OAI22_X1 U2179 ( .A1(n1802), .A2(n2215), .B1(b[21]), .B2(n2215), .ZN(n2214)
         );
  AOI22_X1 U2180 ( .A1(n1805), .A2(n1803), .B1(n1838), .B2(n1803), .ZN(n2215)
         );
  XNOR2_X1 U2181 ( .A(n2219), .B(n1762), .ZN(n714) );
  OAI21_X1 U2182 ( .B1(n1836), .B2(n1792), .A(n2220), .ZN(n2219) );
  OAI22_X1 U2183 ( .A1(n1802), .A2(n2172), .B1(b[22]), .B2(n2172), .ZN(n2220)
         );
  XNOR2_X1 U2184 ( .A(n2222), .B(n1762), .ZN(n713) );
  OAI21_X1 U2185 ( .B1(n1888), .B2(n1792), .A(n2169), .ZN(n2222) );
  XNOR2_X1 U2186 ( .A(a[18]), .B(a[19]), .ZN(n2221) );
  XNOR2_X1 U2187 ( .A(a[19]), .B(n1762), .ZN(n2216) );
  XOR2_X1 U2188 ( .A(a[18]), .B(n1765), .Z(n2217) );
  AOI222_X1 U2189 ( .A1(n2223), .A2(n686), .B1(n1794), .B2(n1745), .C1(n1797), 
        .C2(n1716), .ZN(n711) );
  AOI221_X1 U2190 ( .B1(n1794), .B2(n1649), .C1(n1797), .C2(n1745), .A(n2225), 
        .ZN(n710) );
  OAI22_X1 U2191 ( .A1(n1873), .A2(n1799), .B1(n1775), .B2(n1795), .ZN(n2225)
         );
  OAI22_X1 U2192 ( .A1(n1871), .A2(n1799), .B1(n1876), .B2(n1795), .ZN(n2226)
         );
  AOI221_X1 U2193 ( .B1(n1794), .B2(b[4]), .C1(n1797), .C2(b[3]), .A(n2227), 
        .ZN(n708) );
  OAI22_X1 U2194 ( .A1(n1869), .A2(n1799), .B1(n1874), .B2(n1795), .ZN(n2227)
         );
  AOI221_X1 U2195 ( .B1(n1794), .B2(b[5]), .C1(n1797), .C2(b[4]), .A(n2228), 
        .ZN(n707) );
  OAI22_X1 U2196 ( .A1(n1867), .A2(n1799), .B1(n1872), .B2(n1795), .ZN(n2228)
         );
  AOI221_X1 U2197 ( .B1(n1794), .B2(b[6]), .C1(n1797), .C2(b[5]), .A(n2229), 
        .ZN(n706) );
  OAI22_X1 U2198 ( .A1(n1865), .A2(n1799), .B1(n1870), .B2(n1795), .ZN(n2229)
         );
  AOI221_X1 U2199 ( .B1(n1794), .B2(b[7]), .C1(n1797), .C2(b[6]), .A(n2230), 
        .ZN(n705) );
  OAI22_X1 U2200 ( .A1(n1863), .A2(n1799), .B1(n1868), .B2(n1795), .ZN(n2230)
         );
  AOI221_X1 U2201 ( .B1(n1794), .B2(b[8]), .C1(n1797), .C2(b[7]), .A(n2231), 
        .ZN(n704) );
  OAI22_X1 U2202 ( .A1(n1861), .A2(n1799), .B1(n1866), .B2(n1795), .ZN(n2231)
         );
  AOI221_X1 U2203 ( .B1(n1794), .B2(b[9]), .C1(n1797), .C2(b[8]), .A(n2232), 
        .ZN(n703) );
  OAI22_X1 U2204 ( .A1(n1859), .A2(n1799), .B1(n1864), .B2(n1795), .ZN(n2232)
         );
  AOI221_X1 U2205 ( .B1(n1794), .B2(b[10]), .C1(n1797), .C2(b[9]), .A(n2233), 
        .ZN(n702) );
  OAI22_X1 U2206 ( .A1(n1857), .A2(n1799), .B1(n1862), .B2(n1795), .ZN(n2233)
         );
  AOI221_X1 U2207 ( .B1(n1794), .B2(b[11]), .C1(n1797), .C2(b[10]), .A(n2234), 
        .ZN(n701) );
  OAI22_X1 U2208 ( .A1(n1855), .A2(n1799), .B1(n1860), .B2(n1795), .ZN(n2234)
         );
  AOI221_X1 U2209 ( .B1(n1794), .B2(b[12]), .C1(n1797), .C2(b[11]), .A(n2235), 
        .ZN(n700) );
  OAI22_X1 U2210 ( .A1(n1853), .A2(n1799), .B1(n1858), .B2(n1795), .ZN(n2235)
         );
  AOI221_X1 U2211 ( .B1(n1793), .B2(b[13]), .C1(n1797), .C2(b[12]), .A(n2236), 
        .ZN(n699) );
  OAI22_X1 U2212 ( .A1(n1851), .A2(n1799), .B1(n1856), .B2(n1795), .ZN(n2236)
         );
  AOI221_X1 U2213 ( .B1(n1793), .B2(b[14]), .C1(n1797), .C2(b[13]), .A(n2237), 
        .ZN(n698) );
  OAI22_X1 U2214 ( .A1(n1849), .A2(n1799), .B1(n1854), .B2(n1795), .ZN(n2237)
         );
  AOI221_X1 U2215 ( .B1(n1793), .B2(b[15]), .C1(n1797), .C2(b[14]), .A(n2238), 
        .ZN(n697) );
  OAI22_X1 U2216 ( .A1(n1632), .A2(n1799), .B1(n1852), .B2(n1795), .ZN(n2238)
         );
  AOI221_X1 U2217 ( .B1(n1793), .B2(b[16]), .C1(n1797), .C2(b[15]), .A(n2239), 
        .ZN(n696) );
  OAI22_X1 U2218 ( .A1(n1846), .A2(n1799), .B1(n1850), .B2(n1795), .ZN(n2239)
         );
  AOI221_X1 U2219 ( .B1(n1793), .B2(b[17]), .C1(n1797), .C2(b[16]), .A(n2240), 
        .ZN(n695) );
  OAI22_X1 U2220 ( .A1(n1634), .A2(n1799), .B1(n1848), .B2(n1795), .ZN(n2240)
         );
  AOI221_X1 U2221 ( .B1(n1793), .B2(b[18]), .C1(n1797), .C2(b[17]), .A(n2241), 
        .ZN(n694) );
  OAI22_X1 U2222 ( .A1(n1843), .A2(n1799), .B1(n1847), .B2(n1795), .ZN(n2241)
         );
  AOI221_X1 U2223 ( .B1(n1793), .B2(b[19]), .C1(n1797), .C2(b[18]), .A(n2242), 
        .ZN(n693) );
  OAI22_X1 U2224 ( .A1(n1493), .A2(n1799), .B1(n1845), .B2(n1795), .ZN(n2242)
         );
  AOI221_X1 U2225 ( .B1(n1793), .B2(b[20]), .C1(n1797), .C2(b[19]), .A(n2243), 
        .ZN(n692) );
  OAI22_X1 U2226 ( .A1(n1840), .A2(n1799), .B1(n1844), .B2(n1795), .ZN(n2243)
         );
  AOI221_X1 U2227 ( .B1(n1793), .B2(b[21]), .C1(n1797), .C2(b[20]), .A(n2244), 
        .ZN(n691) );
  OAI22_X1 U2228 ( .A1(n1494), .A2(n1799), .B1(n1842), .B2(n1795), .ZN(n2244)
         );
  OAI22_X1 U2229 ( .A1(n1841), .A2(n1795), .B1(n1839), .B2(n2246), .ZN(n2245)
         );
  AOI22_X1 U2230 ( .A1(n2223), .A2(n2218), .B1(n2247), .B2(n2248), .ZN(n689)
         );
  NAND2_X1 U2231 ( .A1(n2249), .A2(n1839), .ZN(n2248) );
  NAND2_X1 U2232 ( .A1(n2249), .A2(n1795), .ZN(n2247) );
  OAI22_X1 U2233 ( .A1(n1797), .A2(n1794), .B1(b[22]), .B2(n1793), .ZN(n2249)
         );
  XOR2_X1 U2234 ( .A(n641), .B(n1838), .Z(n2218) );
  AOI22_X1 U2235 ( .A1(n2223), .A2(n1888), .B1(n2250), .B2(n2251), .ZN(n688)
         );
  NAND2_X1 U2236 ( .A1(n2246), .A2(n1838), .ZN(n2251) );
  NAND2_X1 U2237 ( .A1(n2246), .A2(n1795), .ZN(n2250) );
  NAND2_X1 U2238 ( .A1(n2253), .A2(n2254), .ZN(n2246) );
  AOI21_X1 U2239 ( .B1(n2223), .B2(n1836), .A(n2252), .ZN(n687) );
  NOR3_X1 U2240 ( .A1(n1800), .A2(a[22]), .A3(n2254), .ZN(n2252) );
  XOR2_X1 U2241 ( .A(a[21]), .B(a[22]), .Z(n2254) );
  NOR2_X1 U2242 ( .A1(n641), .A2(b[22]), .ZN(n1888) );
  AOI22_X1 U2243 ( .A1(n1716), .A2(n1793), .B1(n1716), .B2(n2223), .ZN(n434)
         );
  NOR2_X1 U2244 ( .A1(n2253), .A2(a[22]), .ZN(n2223) );
  AND2_X1 U2245 ( .A1(a[22]), .A2(n1800), .ZN(n2224) );
  XOR2_X1 U2246 ( .A(a[21]), .B(n1763), .Z(n2253) );
  OAI222_X1 U2247 ( .A1(n2256), .A2(n1682), .B1(n2255), .B2(n1796), .C1(n2256), 
        .C2(n1796), .ZN(n150) );
  XNOR2_X1 U2248 ( .A(n2257), .B(n1496), .ZN(n2256) );
  OAI22_X1 U2249 ( .A1(n1600), .A2(n1830), .B1(n1841), .B2(n1733), .ZN(n2258)
         );
  XNOR2_X1 U2250 ( .A(n1482), .B(n2261), .ZN(n2260) );
  OAI22_X1 U2251 ( .A1(n1830), .A2(n1628), .B1(n1842), .B2(n1733), .ZN(n2262)
         );
  OAI222_X1 U2252 ( .A1(n2264), .A2(n2263), .B1(n2263), .B2(n1801), .C1(n2264), 
        .C2(n1801), .ZN(n2259) );
  XNOR2_X1 U2253 ( .A(n1496), .B(n2265), .ZN(n2264) );
  OAI22_X1 U2254 ( .A1(n1830), .A2(n1485), .B1(n1844), .B2(n1733), .ZN(n2266)
         );
  XNOR2_X1 U2255 ( .A(n2269), .B(n1482), .ZN(n2268) );
  AOI221_X1 U2256 ( .B1(n1829), .B2(b[19]), .C1(n1832), .C2(b[18]), .A(n2270), 
        .ZN(n2269) );
  OAI22_X1 U2257 ( .A1(n1830), .A2(n1630), .B1(n1845), .B2(n1733), .ZN(n2270)
         );
  OAI222_X1 U2258 ( .A1(n2272), .A2(n2271), .B1(n2271), .B2(n1476), .C1(n2272), 
        .C2(n1476), .ZN(n2267) );
  XNOR2_X1 U2259 ( .A(n1496), .B(n2273), .ZN(n2272) );
  OAI22_X1 U2260 ( .A1(n1830), .A2(n1495), .B1(n1847), .B2(n1733), .ZN(n2274)
         );
  XNOR2_X1 U2261 ( .A(n1482), .B(n2276), .ZN(n2275) );
  OAI22_X1 U2262 ( .A1(n1830), .A2(n1634), .B1(n1848), .B2(n1733), .ZN(n2277)
         );
  XNOR2_X1 U2263 ( .A(n1496), .B(n2280), .ZN(n2279) );
  OAI22_X1 U2264 ( .A1(n1846), .A2(n1830), .B1(n1850), .B2(n1733), .ZN(n2281)
         );
  XNOR2_X1 U2265 ( .A(n1482), .B(n2284), .ZN(n2283) );
  AOI221_X1 U2266 ( .B1(n1829), .B2(b[15]), .C1(n1832), .C2(b[14]), .A(n2285), 
        .ZN(n2284) );
  OAI22_X1 U2267 ( .A1(n1830), .A2(n1632), .B1(n1852), .B2(n1733), .ZN(n2285)
         );
  OAI222_X1 U2268 ( .A1(n2286), .A2(n2287), .B1(n2286), .B2(n1475), .C1(n1475), 
        .C2(n2287), .ZN(n2282) );
  XNOR2_X1 U2269 ( .A(n2288), .B(n1496), .ZN(n2287) );
  AOI221_X1 U2270 ( .B1(n1829), .B2(b[14]), .C1(n1832), .C2(b[13]), .A(n2289), 
        .ZN(n2288) );
  OAI22_X1 U2271 ( .A1(n1830), .A2(n1849), .B1(n1854), .B2(n1733), .ZN(n2289)
         );
  XNOR2_X1 U2272 ( .A(n1482), .B(n2292), .ZN(n2291) );
  AOI221_X1 U2273 ( .B1(n1829), .B2(b[13]), .C1(n1832), .C2(b[12]), .A(n2293), 
        .ZN(n2292) );
  OAI22_X1 U2274 ( .A1(n1830), .A2(n1851), .B1(n1856), .B2(n1733), .ZN(n2293)
         );
  OAI222_X1 U2275 ( .A1(n2295), .A2(n2296), .B1(n2295), .B2(n1474), .C1(n1474), 
        .C2(n2296), .ZN(n2290) );
  XNOR2_X1 U2276 ( .A(n1496), .B(n2297), .ZN(n2296) );
  AOI221_X1 U2277 ( .B1(n1832), .B2(b[11]), .C1(n675), .C2(n2294), .A(n2298), 
        .ZN(n2297) );
  OAI22_X1 U2278 ( .A1(n1858), .A2(n1733), .B1(n1854), .B2(n1883), .ZN(n2298)
         );
  AOI222_X1 U2279 ( .A1(n2299), .A2(n2300), .B1(n2299), .B2(n527), .C1(n527), 
        .C2(n2300), .ZN(n2295) );
  XNOR2_X1 U2280 ( .A(a[2]), .B(n2301), .ZN(n2300) );
  AOI221_X1 U2281 ( .B1(n1832), .B2(b[10]), .C1(n676), .C2(n2294), .A(n2302), 
        .ZN(n2301) );
  OAI22_X1 U2282 ( .A1(n1856), .A2(n1883), .B1(n1860), .B2(n1733), .ZN(n2302)
         );
  OAI222_X1 U2283 ( .A1(n2303), .A2(n2304), .B1(n2303), .B2(n1817), .C1(n1817), 
        .C2(n2304), .ZN(n2299) );
  XNOR2_X1 U2284 ( .A(n1831), .B(n2305), .ZN(n2304) );
  AOI221_X1 U2285 ( .B1(n1829), .B2(b[10]), .C1(n677), .C2(n2294), .A(n2306), 
        .ZN(n2305) );
  OAI22_X1 U2286 ( .A1(n1860), .A2(n1884), .B1(n1862), .B2(n1733), .ZN(n2306)
         );
  AOI222_X1 U2287 ( .A1(n2307), .A2(n2308), .B1(n2307), .B2(n539), .C1(n539), 
        .C2(n2308), .ZN(n2303) );
  XNOR2_X1 U2288 ( .A(a[2]), .B(n2309), .ZN(n2308) );
  AOI221_X1 U2289 ( .B1(n1829), .B2(b[9]), .C1(n678), .C2(n2294), .A(n2310), 
        .ZN(n2309) );
  OAI22_X1 U2290 ( .A1(n1862), .A2(n1884), .B1(n1864), .B2(n1733), .ZN(n2310)
         );
  OAI222_X1 U2291 ( .A1(n2311), .A2(n2312), .B1(n2311), .B2(n1822), .C1(n1822), 
        .C2(n2312), .ZN(n2307) );
  XNOR2_X1 U2292 ( .A(n1831), .B(n2313), .ZN(n2312) );
  AOI221_X1 U2293 ( .B1(n1829), .B2(b[8]), .C1(n679), .C2(n2294), .A(n2314), 
        .ZN(n2313) );
  OAI22_X1 U2294 ( .A1(n1864), .A2(n1884), .B1(n1866), .B2(n1733), .ZN(n2314)
         );
  XNOR2_X1 U2295 ( .A(a[2]), .B(n2317), .ZN(n2316) );
  AOI221_X1 U2296 ( .B1(n1829), .B2(b[7]), .C1(n680), .C2(n2294), .A(n2318), 
        .ZN(n2317) );
  OAI22_X1 U2297 ( .A1(n1866), .A2(n1884), .B1(n1868), .B2(n1733), .ZN(n2318)
         );
  OAI222_X1 U2298 ( .A1(n2319), .A2(n2320), .B1(n2319), .B2(n1823), .C1(n1823), 
        .C2(n2320), .ZN(n2315) );
  XNOR2_X1 U2299 ( .A(n1831), .B(n2321), .ZN(n2320) );
  AOI221_X1 U2300 ( .B1(n1829), .B2(b[6]), .C1(n681), .C2(n2294), .A(n2322), 
        .ZN(n2321) );
  OAI22_X1 U2301 ( .A1(n1868), .A2(n1884), .B1(n1870), .B2(n1733), .ZN(n2322)
         );
  AOI222_X1 U2302 ( .A1(n2323), .A2(n2324), .B1(n2323), .B2(n557), .C1(n557), 
        .C2(n2324), .ZN(n2319) );
  XNOR2_X1 U2303 ( .A(a[2]), .B(n2325), .ZN(n2324) );
  AOI221_X1 U2304 ( .B1(n1829), .B2(b[5]), .C1(n682), .C2(n2294), .A(n2326), 
        .ZN(n2325) );
  OAI22_X1 U2305 ( .A1(n1870), .A2(n1884), .B1(n1872), .B2(n1733), .ZN(n2326)
         );
  OAI222_X1 U2306 ( .A1(n2327), .A2(n2328), .B1(n2327), .B2(n1826), .C1(n1826), 
        .C2(n2328), .ZN(n2323) );
  XNOR2_X1 U2307 ( .A(n1831), .B(n2329), .ZN(n2328) );
  AOI221_X1 U2308 ( .B1(n1829), .B2(b[4]), .C1(n683), .C2(n2294), .A(n2330), 
        .ZN(n2329) );
  OAI22_X1 U2309 ( .A1(n1872), .A2(n1884), .B1(n1874), .B2(n1733), .ZN(n2330)
         );
  XNOR2_X1 U2310 ( .A(a[2]), .B(n2333), .ZN(n2332) );
  AOI221_X1 U2311 ( .B1(n1829), .B2(b[3]), .C1(n684), .C2(n2294), .A(n2334), 
        .ZN(n2333) );
  OAI22_X1 U2312 ( .A1(n1874), .A2(n1884), .B1(n1876), .B2(n1733), .ZN(n2334)
         );
  AND4_X1 U2313 ( .A1(a[2]), .A2(n1776), .A3(n2336), .A4(n2337), .ZN(n2331) );
  AOI222_X1 U2314 ( .A1(n685), .A2(n2294), .B1(n1832), .B2(n1602), .C1(n1829), 
        .C2(n1649), .ZN(n2337) );
  AOI22_X1 U2315 ( .A1(n1829), .A2(n1602), .B1(n686), .B2(n2294), .ZN(n2336)
         );
  XNOR2_X1 U2316 ( .A(n1833), .B(n1831), .ZN(n2335) );
endmodule


module FPMultiplier ( clk, a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input clk;
  wire   N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, N3, add_0_root_sub_1_root_sub_23_A_0_,
         add_0_root_sub_1_root_sub_23_A_1_, add_0_root_sub_1_root_sub_23_A_2_,
         add_0_root_sub_1_root_sub_23_A_3_, add_0_root_sub_1_root_sub_23_A_4_,
         add_0_root_sub_1_root_sub_23_A_5_, add_0_root_sub_1_root_sub_23_A_6_,
         add_0_root_sub_1_root_sub_23_A_7_, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23;
  wire   [31:0] a_reg;
  wire   [31:0] b_reg;
  wire   [46:23] tempMantisa;
  wire   [7:2] add_0_root_sub_1_root_sub_23_carry;

  DFF_X1 a_reg_reg_31_ ( .D(a[31]), .CK(clk), .Q(a_reg[31]) );
  DFF_X1 a_reg_reg_30_ ( .D(a[30]), .CK(clk), .Q(a_reg[30]) );
  DFF_X1 a_reg_reg_29_ ( .D(a[29]), .CK(clk), .Q(a_reg[29]) );
  DFF_X1 a_reg_reg_28_ ( .D(a[28]), .CK(clk), .Q(a_reg[28]) );
  DFF_X1 a_reg_reg_27_ ( .D(a[27]), .CK(clk), .Q(a_reg[27]) );
  DFF_X1 a_reg_reg_26_ ( .D(a[26]), .CK(clk), .Q(a_reg[26]) );
  DFF_X1 a_reg_reg_25_ ( .D(a[25]), .CK(clk), .Q(a_reg[25]) );
  DFF_X1 a_reg_reg_24_ ( .D(a[24]), .CK(clk), .Q(a_reg[24]) );
  DFF_X1 a_reg_reg_23_ ( .D(a[23]), .CK(clk), .Q(a_reg[23]) );
  DFF_X1 a_reg_reg_22_ ( .D(a[22]), .CK(clk), .Q(a_reg[22]) );
  DFF_X1 a_reg_reg_21_ ( .D(a[21]), .CK(clk), .Q(a_reg[21]) );
  DFF_X1 a_reg_reg_20_ ( .D(a[20]), .CK(clk), .Q(a_reg[20]) );
  DFF_X1 a_reg_reg_19_ ( .D(a[19]), .CK(clk), .Q(a_reg[19]) );
  DFF_X1 a_reg_reg_18_ ( .D(a[18]), .CK(clk), .Q(a_reg[18]) );
  DFF_X1 a_reg_reg_17_ ( .D(a[17]), .CK(clk), .Q(a_reg[17]) );
  DFF_X1 a_reg_reg_16_ ( .D(a[16]), .CK(clk), .Q(a_reg[16]) );
  DFF_X1 a_reg_reg_15_ ( .D(a[15]), .CK(clk), .Q(a_reg[15]) );
  DFF_X1 a_reg_reg_14_ ( .D(a[14]), .CK(clk), .Q(a_reg[14]) );
  DFF_X1 a_reg_reg_13_ ( .D(a[13]), .CK(clk), .Q(a_reg[13]) );
  DFF_X1 a_reg_reg_12_ ( .D(a[12]), .CK(clk), .Q(a_reg[12]) );
  DFF_X1 a_reg_reg_11_ ( .D(a[11]), .CK(clk), .Q(a_reg[11]) );
  DFF_X1 a_reg_reg_10_ ( .D(a[10]), .CK(clk), .Q(a_reg[10]) );
  DFF_X1 a_reg_reg_9_ ( .D(a[9]), .CK(clk), .Q(a_reg[9]) );
  DFF_X1 a_reg_reg_8_ ( .D(a[8]), .CK(clk), .Q(a_reg[8]) );
  DFF_X1 a_reg_reg_7_ ( .D(a[7]), .CK(clk), .Q(a_reg[7]) );
  DFF_X1 a_reg_reg_6_ ( .D(a[6]), .CK(clk), .Q(a_reg[6]) );
  DFF_X1 a_reg_reg_5_ ( .D(a[5]), .CK(clk), .Q(a_reg[5]), .QN(n72) );
  DFF_X1 a_reg_reg_4_ ( .D(a[4]), .CK(clk), .Q(a_reg[4]) );
  DFF_X1 a_reg_reg_3_ ( .D(a[3]), .CK(clk), .Q(a_reg[3]) );
  DFF_X1 a_reg_reg_1_ ( .D(a[1]), .CK(clk), .Q(a_reg[1]) );
  DFF_X1 a_reg_reg_0_ ( .D(a[0]), .CK(clk), .Q(a_reg[0]) );
  DFF_X1 b_reg_reg_31_ ( .D(b[31]), .CK(clk), .Q(b_reg[31]) );
  DFF_X1 result_reg_31_ ( .D(N81), .CK(clk), .Q(result[31]) );
  DFF_X1 b_reg_reg_30_ ( .D(b[30]), .CK(clk), .Q(b_reg[30]) );
  DFF_X1 b_reg_reg_29_ ( .D(b[29]), .CK(clk), .Q(b_reg[29]) );
  DFF_X1 b_reg_reg_28_ ( .D(b[28]), .CK(clk), .Q(b_reg[28]) );
  DFF_X1 b_reg_reg_27_ ( .D(b[27]), .CK(clk), .Q(b_reg[27]) );
  DFF_X1 b_reg_reg_26_ ( .D(b[26]), .CK(clk), .Q(b_reg[26]) );
  DFF_X1 b_reg_reg_25_ ( .D(b[25]), .CK(clk), .Q(b_reg[25]) );
  DFF_X1 b_reg_reg_24_ ( .D(b[24]), .CK(clk), .Q(b_reg[24]) );
  DFF_X1 b_reg_reg_23_ ( .D(b[23]), .CK(clk), .Q(b_reg[23]) );
  DFF_X1 b_reg_reg_22_ ( .D(b[22]), .CK(clk), .Q(b_reg[22]) );
  DFF_X1 b_reg_reg_21_ ( .D(b[21]), .CK(clk), .Q(b_reg[21]) );
  DFF_X1 b_reg_reg_20_ ( .D(b[20]), .CK(clk), .Q(b_reg[20]) );
  DFF_X1 b_reg_reg_19_ ( .D(b[19]), .CK(clk), .Q(b_reg[19]) );
  DFF_X1 b_reg_reg_18_ ( .D(b[18]), .CK(clk), .Q(b_reg[18]) );
  DFF_X1 b_reg_reg_17_ ( .D(b[17]), .CK(clk), .Q(b_reg[17]) );
  DFF_X1 b_reg_reg_16_ ( .D(b[16]), .CK(clk), .Q(b_reg[16]) );
  DFF_X1 b_reg_reg_15_ ( .D(b[15]), .CK(clk), .Q(b_reg[15]) );
  DFF_X1 b_reg_reg_14_ ( .D(b[14]), .CK(clk), .Q(b_reg[14]) );
  DFF_X1 b_reg_reg_13_ ( .D(b[13]), .CK(clk), .Q(b_reg[13]) );
  DFF_X1 b_reg_reg_12_ ( .D(b[12]), .CK(clk), .Q(b_reg[12]) );
  DFF_X1 b_reg_reg_11_ ( .D(b[11]), .CK(clk), .Q(b_reg[11]) );
  DFF_X1 b_reg_reg_10_ ( .D(b[10]), .CK(clk), .Q(b_reg[10]) );
  DFF_X1 b_reg_reg_9_ ( .D(b[9]), .CK(clk), .Q(b_reg[9]) );
  DFF_X1 b_reg_reg_8_ ( .D(b[8]), .CK(clk), .Q(b_reg[8]) );
  DFF_X1 b_reg_reg_7_ ( .D(b[7]), .CK(clk), .Q(b_reg[7]) );
  DFF_X1 b_reg_reg_6_ ( .D(b[6]), .CK(clk), .Q(b_reg[6]) );
  DFF_X1 b_reg_reg_5_ ( .D(b[5]), .CK(clk), .Q(b_reg[5]) );
  DFF_X1 b_reg_reg_4_ ( .D(b[4]), .CK(clk), .Q(b_reg[4]) );
  DFF_X1 b_reg_reg_0_ ( .D(b[0]), .CK(clk), .Q(b_reg[0]), .QN(n54) );
  DFF_X1 result_reg_23_ ( .D(N33), .CK(clk), .Q(result[23]) );
  DFF_X1 result_reg_24_ ( .D(N32), .CK(clk), .Q(result[24]) );
  DFF_X1 result_reg_25_ ( .D(N31), .CK(clk), .Q(result[25]) );
  DFF_X1 result_reg_26_ ( .D(N30), .CK(clk), .Q(result[26]) );
  DFF_X1 result_reg_27_ ( .D(N29), .CK(clk), .Q(result[27]) );
  DFF_X1 result_reg_28_ ( .D(N28), .CK(clk), .Q(result[28]) );
  DFF_X1 result_reg_29_ ( .D(N27), .CK(clk), .Q(result[29]) );
  DFF_X1 result_reg_0_ ( .D(N80), .CK(clk), .Q(result[0]) );
  DFF_X1 result_reg_1_ ( .D(N79), .CK(clk), .Q(result[1]) );
  DFF_X1 result_reg_2_ ( .D(N78), .CK(clk), .Q(result[2]) );
  DFF_X1 result_reg_3_ ( .D(N77), .CK(clk), .Q(result[3]) );
  DFF_X1 result_reg_4_ ( .D(N76), .CK(clk), .Q(result[4]) );
  DFF_X1 result_reg_5_ ( .D(N75), .CK(clk), .Q(result[5]) );
  DFF_X1 result_reg_6_ ( .D(N74), .CK(clk), .Q(result[6]) );
  DFF_X1 result_reg_7_ ( .D(N73), .CK(clk), .Q(result[7]) );
  DFF_X1 result_reg_8_ ( .D(N72), .CK(clk), .Q(result[8]) );
  DFF_X1 result_reg_9_ ( .D(N71), .CK(clk), .Q(result[9]) );
  DFF_X1 result_reg_10_ ( .D(N70), .CK(clk), .Q(result[10]) );
  DFF_X1 result_reg_11_ ( .D(N69), .CK(clk), .Q(result[11]) );
  DFF_X1 result_reg_12_ ( .D(N68), .CK(clk), .Q(result[12]) );
  DFF_X1 result_reg_13_ ( .D(N67), .CK(clk), .Q(result[13]) );
  DFF_X1 result_reg_14_ ( .D(N66), .CK(clk), .Q(result[14]) );
  DFF_X1 result_reg_15_ ( .D(N65), .CK(clk), .Q(result[15]) );
  DFF_X1 result_reg_16_ ( .D(N64), .CK(clk), .Q(result[16]) );
  DFF_X1 result_reg_17_ ( .D(N63), .CK(clk), .Q(result[17]) );
  DFF_X1 result_reg_18_ ( .D(N62), .CK(clk), .Q(result[18]) );
  DFF_X1 result_reg_19_ ( .D(N61), .CK(clk), .Q(result[19]) );
  DFF_X1 result_reg_20_ ( .D(N60), .CK(clk), .Q(result[20]) );
  DFF_X1 result_reg_21_ ( .D(N59), .CK(clk), .Q(result[21]) );
  DFF_X1 result_reg_22_ ( .D(N58), .CK(clk), .Q(result[22]) );
  XOR2_X1 U82 ( .A(b_reg[31]), .B(a_reg[31]), .Z(N81) );
  FPMultiplier_DW01_add_1 add_2_root_sub_1_root_sub_23 ( .A(b_reg[30:23]), .B(
        a_reg[30:23]), .CI(1'b0), .SUM({add_0_root_sub_1_root_sub_23_A_7_, 
        add_0_root_sub_1_root_sub_23_A_6_, add_0_root_sub_1_root_sub_23_A_5_, 
        add_0_root_sub_1_root_sub_23_A_4_, add_0_root_sub_1_root_sub_23_A_3_, 
        add_0_root_sub_1_root_sub_23_A_2_, add_0_root_sub_1_root_sub_23_A_1_, 
        add_0_root_sub_1_root_sub_23_A_0_}) );
  FPMultiplier_DW_mult_uns_0 mult_17 ( .a({1'b1, a_reg[22:3], n61, a_reg[1:0]}), .b({1'b1, b_reg[22:0]}), .product({N3, tempMantisa, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23}) );
  FA_X1 add_0_root_sub_1_root_sub_23_U1_1 ( .A(n68), .B(
        add_0_root_sub_1_root_sub_23_A_1_), .CI(n71), .CO(
        add_0_root_sub_1_root_sub_23_carry[2]), .S(N19) );
  DFF_X1 b_reg_reg_2_ ( .D(b[2]), .CK(clk), .Q(b_reg[2]) );
  DFF_X1 result_reg_30_ ( .D(N26), .CK(clk), .Q(result[30]) );
  DFF_X2 b_reg_reg_3_ ( .D(b[3]), .CK(clk), .Q(b_reg[3]) );
  DFF_X1 a_reg_reg_2_ ( .D(a[2]), .CK(clk), .Q(a_reg[2]) );
  DFF_X1 b_reg_reg_1_ ( .D(b[1]), .CK(clk), .Q(b_reg[1]), .QN(n56) );
  FA_X1 add_0_root_sub_1_root_sub_23_U1_4 ( .A(
        add_0_root_sub_1_root_sub_23_A_4_), .B(1'b0), .CI(
        add_0_root_sub_1_root_sub_23_carry[4]), .CO(
        add_0_root_sub_1_root_sub_23_carry[5]), .S(N22) );
  INV_X2 U83 ( .A(n65), .ZN(add_0_root_sub_1_root_sub_23_carry[7]) );
  INV_X2 U84 ( .A(n66), .ZN(add_0_root_sub_1_root_sub_23_carry[6]) );
  INV_X2 U85 ( .A(n66), .ZN(n63) );
  INV_X2 U86 ( .A(n64), .ZN(add_0_root_sub_1_root_sub_23_carry[4]) );
  INV_X2 U87 ( .A(n58), .ZN(add_0_root_sub_1_root_sub_23_carry[3]) );
  AND2_X1 U88 ( .A1(n69), .A2(n76), .ZN(N33) );
  BUF_X2 U89 ( .A(a_reg[2]), .Z(n61) );
  CLKBUF_X1 U90 ( .A(add_0_root_sub_1_root_sub_23_carry[2]), .Z(n53) );
  INV_X1 U91 ( .A(n54), .ZN(n55) );
  INV_X1 U92 ( .A(n56), .ZN(n57) );
  XOR2_X1 U93 ( .A(n53), .B(add_0_root_sub_1_root_sub_23_A_2_), .Z(N20) );
  NAND2_X1 U94 ( .A1(add_0_root_sub_1_root_sub_23_carry[2]), .A2(
        add_0_root_sub_1_root_sub_23_A_2_), .ZN(n58) );
  INV_X1 U95 ( .A(n67), .ZN(n59) );
  CLKBUF_X1 U96 ( .A(add_0_root_sub_1_root_sub_23_carry[5]), .Z(n60) );
  CLKBUF_X1 U97 ( .A(add_0_root_sub_1_root_sub_23_carry[3]), .Z(n62) );
  XOR2_X1 U98 ( .A(n62), .B(add_0_root_sub_1_root_sub_23_A_3_), .Z(N21) );
  NAND2_X1 U99 ( .A1(add_0_root_sub_1_root_sub_23_carry[3]), .A2(
        add_0_root_sub_1_root_sub_23_A_3_), .ZN(n64) );
  XOR2_X1 U100 ( .A(n63), .B(add_0_root_sub_1_root_sub_23_A_6_), .Z(N24) );
  NAND2_X1 U101 ( .A1(add_0_root_sub_1_root_sub_23_carry[6]), .A2(
        add_0_root_sub_1_root_sub_23_A_6_), .ZN(n65) );
  XOR2_X1 U102 ( .A(n60), .B(add_0_root_sub_1_root_sub_23_A_5_), .Z(N23) );
  NAND2_X1 U103 ( .A1(add_0_root_sub_1_root_sub_23_carry[5]), .A2(
        add_0_root_sub_1_root_sub_23_A_5_), .ZN(n66) );
  CLKBUF_X1 U104 ( .A(n71), .Z(n67) );
  OAI22_X1 U105 ( .A1(n74), .A2(n89), .B1(n75), .B2(n90), .ZN(N70) );
  OAI22_X1 U106 ( .A1(n74), .A2(n93), .B1(n75), .B2(n94), .ZN(N74) );
  OAI22_X1 U107 ( .A1(n74), .A2(n95), .B1(n75), .B2(n96), .ZN(N76) );
  OAI22_X1 U108 ( .A1(n74), .A2(n97), .B1(n75), .B2(n98), .ZN(N78) );
  OAI22_X1 U109 ( .A1(n30), .A2(n86), .B1(n31), .B2(n87), .ZN(N67) );
  OAI22_X1 U110 ( .A1(n30), .A2(n94), .B1(n31), .B2(n95), .ZN(N75) );
  OAI22_X1 U111 ( .A1(n30), .A2(n96), .B1(n31), .B2(n97), .ZN(N77) );
  OAI22_X1 U112 ( .A1(n74), .A2(n79), .B1(n75), .B2(n80), .ZN(N60) );
  OAI22_X1 U113 ( .A1(n74), .A2(n81), .B1(n75), .B2(n82), .ZN(N62) );
  OAI22_X1 U114 ( .A1(n74), .A2(n83), .B1(n75), .B2(n84), .ZN(N64) );
  OAI22_X1 U115 ( .A1(n74), .A2(n85), .B1(n75), .B2(n86), .ZN(N66) );
  OAI22_X1 U116 ( .A1(n74), .A2(n87), .B1(n75), .B2(n88), .ZN(N68) );
  OAI22_X1 U117 ( .A1(n74), .A2(n91), .B1(n75), .B2(n92), .ZN(N72) );
  OAI22_X1 U118 ( .A1(n74), .A2(n99), .B1(n75), .B2(n100), .ZN(N80) );
  INV_X1 U119 ( .A(tempMantisa[23]), .ZN(n100) );
  OAI22_X1 U120 ( .A1(n30), .A2(n78), .B1(n31), .B2(n79), .ZN(N59) );
  OAI22_X1 U121 ( .A1(n30), .A2(n80), .B1(n31), .B2(n81), .ZN(N61) );
  OAI22_X1 U122 ( .A1(n30), .A2(n82), .B1(n31), .B2(n83), .ZN(N63) );
  OAI22_X1 U123 ( .A1(n30), .A2(n84), .B1(n31), .B2(n85), .ZN(N65) );
  OAI22_X1 U124 ( .A1(n30), .A2(n88), .B1(n31), .B2(n89), .ZN(N69) );
  OAI22_X1 U125 ( .A1(n30), .A2(n90), .B1(n31), .B2(n91), .ZN(N71) );
  OAI22_X1 U126 ( .A1(n30), .A2(n92), .B1(n31), .B2(n93), .ZN(N73) );
  OAI22_X1 U127 ( .A1(n30), .A2(n98), .B1(n31), .B2(n99), .ZN(N79) );
  INV_X1 U128 ( .A(tempMantisa[45]), .ZN(n78) );
  INV_X1 U129 ( .A(tempMantisa[43]), .ZN(n80) );
  INV_X1 U130 ( .A(tempMantisa[41]), .ZN(n82) );
  INV_X1 U131 ( .A(tempMantisa[39]), .ZN(n84) );
  AND2_X1 U132 ( .A1(N19), .A2(n76), .ZN(N32) );
  INV_X1 U133 ( .A(tempMantisa[37]), .ZN(n86) );
  INV_X1 U134 ( .A(tempMantisa[36]), .ZN(n87) );
  INV_X1 U135 ( .A(tempMantisa[34]), .ZN(n89) );
  INV_X1 U136 ( .A(tempMantisa[33]), .ZN(n90) );
  INV_X1 U137 ( .A(tempMantisa[30]), .ZN(n93) );
  INV_X1 U138 ( .A(tempMantisa[29]), .ZN(n94) );
  INV_X1 U139 ( .A(tempMantisa[27]), .ZN(n96) );
  INV_X1 U140 ( .A(tempMantisa[26]), .ZN(n97) );
  INV_X1 U141 ( .A(tempMantisa[25]), .ZN(n98) );
  INV_X1 U142 ( .A(tempMantisa[28]), .ZN(n95) );
  INV_X1 U143 ( .A(n32), .ZN(n76) );
  OAI22_X1 U144 ( .A1(n74), .A2(n77), .B1(n75), .B2(n78), .ZN(N58) );
  INV_X1 U145 ( .A(tempMantisa[46]), .ZN(n77) );
  AND2_X1 U146 ( .A1(n70), .A2(add_0_root_sub_1_root_sub_23_A_0_), .ZN(n68) );
  INV_X1 U147 ( .A(tempMantisa[44]), .ZN(n79) );
  INV_X1 U148 ( .A(tempMantisa[40]), .ZN(n83) );
  INV_X1 U149 ( .A(tempMantisa[38]), .ZN(n85) );
  INV_X1 U150 ( .A(tempMantisa[42]), .ZN(n81) );
  AND2_X1 U151 ( .A1(N24), .A2(n76), .ZN(N27) );
  AND2_X1 U152 ( .A1(N20), .A2(n76), .ZN(N31) );
  XOR2_X1 U153 ( .A(n59), .B(add_0_root_sub_1_root_sub_23_A_0_), .Z(n69) );
  AND2_X1 U154 ( .A1(N23), .A2(n76), .ZN(N28) );
  AND2_X1 U155 ( .A1(N22), .A2(n76), .ZN(N29) );
  AND2_X1 U156 ( .A1(N21), .A2(n76), .ZN(N30) );
  INV_X1 U157 ( .A(tempMantisa[35]), .ZN(n88) );
  INV_X1 U158 ( .A(tempMantisa[32]), .ZN(n91) );
  INV_X1 U159 ( .A(tempMantisa[31]), .ZN(n92) );
  INV_X1 U160 ( .A(tempMantisa[24]), .ZN(n99) );
  OAI22_X1 U161 ( .A1(n33), .A2(n34), .B1(n35), .B2(n36), .ZN(n32) );
  NAND4_X1 U162 ( .A1(n41), .A2(n42), .A3(n43), .A4(n44), .ZN(n35) );
  NAND4_X1 U163 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .ZN(n36) );
  NAND4_X1 U164 ( .A1(n49), .A2(n50), .A3(n51), .A4(n52), .ZN(n33) );
  XNOR2_X1 U165 ( .A(add_0_root_sub_1_root_sub_23_carry[7]), .B(
        add_0_root_sub_1_root_sub_23_A_7_), .ZN(N25) );
  NOR4_X1 U166 ( .A1(b_reg[9]), .A2(b_reg[8]), .A3(b_reg[7]), .A4(b_reg[6]), 
        .ZN(n52) );
  NOR4_X1 U167 ( .A1(b_reg[19]), .A2(b_reg[18]), .A3(b_reg[17]), .A4(b_reg[16]), .ZN(n47) );
  NOR4_X1 U168 ( .A1(b_reg[5]), .A2(b_reg[4]), .A3(b_reg[3]), .A4(b_reg[30]), 
        .ZN(n51) );
  NOR4_X1 U169 ( .A1(a_reg[22]), .A2(a_reg[21]), .A3(a_reg[20]), .A4(a_reg[1]), 
        .ZN(n40) );
  NOR4_X1 U170 ( .A1(a_reg[9]), .A2(a_reg[8]), .A3(a_reg[7]), .A4(a_reg[6]), 
        .ZN(n44) );
  NOR4_X1 U171 ( .A1(a_reg[19]), .A2(a_reg[18]), .A3(a_reg[17]), .A4(a_reg[16]), .ZN(n39) );
  NOR4_X1 U172 ( .A1(a_reg[15]), .A2(a_reg[14]), .A3(a_reg[13]), .A4(a_reg[12]), .ZN(n38) );
  NOR4_X1 U173 ( .A1(b_reg[26]), .A2(b_reg[25]), .A3(b_reg[24]), .A4(b_reg[23]), .ZN(n49) );
  NOR4_X1 U174 ( .A1(a_reg[26]), .A2(a_reg[25]), .A3(a_reg[24]), .A4(a_reg[23]), .ZN(n41) );
  NOR3_X1 U175 ( .A1(a_reg[0]), .A2(a_reg[11]), .A3(a_reg[10]), .ZN(n37) );
  NAND4_X1 U176 ( .A1(n45), .A2(n46), .A3(n47), .A4(n48), .ZN(n34) );
  NOR3_X1 U177 ( .A1(n55), .A2(b_reg[11]), .A3(b_reg[10]), .ZN(n45) );
  NOR4_X1 U178 ( .A1(b_reg[15]), .A2(b_reg[14]), .A3(b_reg[13]), .A4(b_reg[12]), .ZN(n46) );
  INV_X1 U179 ( .A(N3), .ZN(n70) );
  INV_X1 U180 ( .A(n70), .ZN(n71) );
  INV_X1 U181 ( .A(n72), .ZN(n73) );
  AND2_X1 U182 ( .A1(N25), .A2(n76), .ZN(N26) );
  NOR4_X1 U183 ( .A1(b_reg[22]), .A2(b_reg[21]), .A3(b_reg[20]), .A4(n57), 
        .ZN(n48) );
  NOR4_X1 U184 ( .A1(n73), .A2(a_reg[4]), .A3(a_reg[3]), .A4(a_reg[30]), .ZN(
        n43) );
  NOR4_X1 U185 ( .A1(b_reg[2]), .A2(b_reg[29]), .A3(b_reg[28]), .A4(b_reg[27]), 
        .ZN(n50) );
  NOR4_X1 U186 ( .A1(n61), .A2(a_reg[29]), .A3(a_reg[28]), .A4(a_reg[27]), 
        .ZN(n42) );
  NAND2_X1 U187 ( .A1(n67), .A2(n76), .ZN(n30) );
  NAND2_X1 U188 ( .A1(n67), .A2(n76), .ZN(n74) );
  OR2_X1 U189 ( .A1(n32), .A2(n67), .ZN(n31) );
  OR2_X1 U190 ( .A1(n32), .A2(n71), .ZN(n75) );
endmodule

