module TopModule (
    input wire clk,
    input wire iclk,
    input wire [31:0] a,
    input wire [31:0] b,
    input  wire reset ,
    input wire resetReg,
    output wire [63:0] result
);
wire [31:0] mulA;
wire [31:0] mulB;
wire [63:0] mulResult;

register #(.N(64)) R0(.clk(clk),.reset(resetReg),.reg_in({a,b}),.reg_out({mulA,mulB}));
//register #(.N(32)) R1(.clk(clk),.reset(resetReg),.reg_in(b),.reg_out(mulB));


boothMultiplier M0(.a(mulA),.b(mulB),.reset(reset),.clk(iclk),.result(mulResult));

register #(.N(64)) R2(.clk(clk),.reset(resetReg),.reg_in(mulResult),.reg_out(result));
    
endmodule

// booth multiplier top module
