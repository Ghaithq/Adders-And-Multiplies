
module register_N32_0 ( clk, reset, reg_in, reg_out );
  input [31:0] reg_in;
  output [31:0] reg_out;
  input clk, reset;
  wire   n33, n34, n35, n36;

  SDFF_X1 reg_out_reg_31_ ( .D(1'b0), .SI(n33), .SE(reg_in[31]), .CK(clk), .Q(
        reg_out[31]) );
  SDFF_X1 reg_out_reg_30_ ( .D(1'b0), .SI(n33), .SE(reg_in[30]), .CK(clk), .Q(
        reg_out[30]) );
  SDFF_X1 reg_out_reg_29_ ( .D(1'b0), .SI(n33), .SE(reg_in[29]), .CK(clk), .Q(
        reg_out[29]) );
  SDFF_X1 reg_out_reg_28_ ( .D(1'b0), .SI(n33), .SE(reg_in[28]), .CK(clk), .Q(
        reg_out[28]) );
  SDFF_X1 reg_out_reg_27_ ( .D(1'b0), .SI(n33), .SE(reg_in[27]), .CK(clk), .Q(
        reg_out[27]) );
  SDFF_X1 reg_out_reg_26_ ( .D(1'b0), .SI(n33), .SE(reg_in[26]), .CK(clk), .Q(
        reg_out[26]) );
  SDFF_X1 reg_out_reg_25_ ( .D(1'b0), .SI(n33), .SE(reg_in[25]), .CK(clk), .Q(
        reg_out[25]) );
  SDFF_X1 reg_out_reg_24_ ( .D(1'b0), .SI(n33), .SE(reg_in[24]), .CK(clk), .Q(
        reg_out[24]) );
  SDFF_X1 reg_out_reg_23_ ( .D(1'b0), .SI(n33), .SE(reg_in[23]), .CK(clk), .Q(
        reg_out[23]) );
  SDFF_X1 reg_out_reg_22_ ( .D(1'b0), .SI(n33), .SE(reg_in[22]), .CK(clk), .Q(
        reg_out[22]) );
  SDFF_X1 reg_out_reg_21_ ( .D(1'b0), .SI(n33), .SE(reg_in[21]), .CK(clk), .Q(
        reg_out[21]) );
  SDFF_X1 reg_out_reg_20_ ( .D(1'b0), .SI(n34), .SE(reg_in[20]), .CK(clk), .Q(
        reg_out[20]) );
  SDFF_X1 reg_out_reg_19_ ( .D(1'b0), .SI(n34), .SE(reg_in[19]), .CK(clk), .Q(
        reg_out[19]) );
  SDFF_X1 reg_out_reg_18_ ( .D(1'b0), .SI(n34), .SE(reg_in[18]), .CK(clk), .Q(
        reg_out[18]) );
  SDFF_X1 reg_out_reg_17_ ( .D(1'b0), .SI(n34), .SE(reg_in[17]), .CK(clk), .Q(
        reg_out[17]) );
  SDFF_X1 reg_out_reg_16_ ( .D(1'b0), .SI(n34), .SE(reg_in[16]), .CK(clk), .Q(
        reg_out[16]) );
  SDFF_X1 reg_out_reg_15_ ( .D(1'b0), .SI(n34), .SE(reg_in[15]), .CK(clk), .Q(
        reg_out[15]) );
  SDFF_X1 reg_out_reg_14_ ( .D(1'b0), .SI(n34), .SE(reg_in[14]), .CK(clk), .Q(
        reg_out[14]) );
  SDFF_X1 reg_out_reg_13_ ( .D(1'b0), .SI(n34), .SE(reg_in[13]), .CK(clk), .Q(
        reg_out[13]) );
  SDFF_X1 reg_out_reg_12_ ( .D(1'b0), .SI(n34), .SE(reg_in[12]), .CK(clk), .Q(
        reg_out[12]) );
  SDFF_X1 reg_out_reg_11_ ( .D(1'b0), .SI(n34), .SE(reg_in[11]), .CK(clk), .Q(
        reg_out[11]) );
  SDFF_X1 reg_out_reg_10_ ( .D(1'b0), .SI(n34), .SE(reg_in[10]), .CK(clk), .Q(
        reg_out[10]) );
  SDFF_X1 reg_out_reg_9_ ( .D(1'b0), .SI(n35), .SE(reg_in[9]), .CK(clk), .Q(
        reg_out[9]) );
  SDFF_X1 reg_out_reg_8_ ( .D(1'b0), .SI(n35), .SE(reg_in[8]), .CK(clk), .Q(
        reg_out[8]) );
  SDFF_X1 reg_out_reg_7_ ( .D(1'b0), .SI(n35), .SE(reg_in[7]), .CK(clk), .Q(
        reg_out[7]) );
  SDFF_X1 reg_out_reg_6_ ( .D(1'b0), .SI(n35), .SE(reg_in[6]), .CK(clk), .Q(
        reg_out[6]) );
  SDFF_X1 reg_out_reg_5_ ( .D(1'b0), .SI(n35), .SE(reg_in[5]), .CK(clk), .Q(
        reg_out[5]) );
  SDFF_X1 reg_out_reg_4_ ( .D(1'b0), .SI(n35), .SE(reg_in[4]), .CK(clk), .Q(
        reg_out[4]) );
  SDFF_X1 reg_out_reg_3_ ( .D(1'b0), .SI(n35), .SE(reg_in[3]), .CK(clk), .Q(
        reg_out[3]) );
  SDFF_X1 reg_out_reg_2_ ( .D(1'b0), .SI(n35), .SE(reg_in[2]), .CK(clk), .Q(
        reg_out[2]) );
  SDFF_X1 reg_out_reg_1_ ( .D(1'b0), .SI(n35), .SE(reg_in[1]), .CK(clk), .Q(
        reg_out[1]) );
  SDFF_X1 reg_out_reg_0_ ( .D(1'b0), .SI(n35), .SE(reg_in[0]), .CK(clk), .Q(
        reg_out[0]) );
  BUF_X1 U35 ( .A(n36), .Z(n34) );
  BUF_X1 U36 ( .A(n36), .Z(n35) );
  INV_X1 U37 ( .A(reset), .ZN(n36) );
  BUF_X1 U38 ( .A(n36), .Z(n33) );
endmodule


module register_N32_1 ( clk, reset, reg_in, reg_out );
  input [31:0] reg_in;
  output [31:0] reg_out;
  input clk, reset;
  wire   n33, n34, n35, n36;

  SDFF_X1 reg_out_reg_31_ ( .D(1'b0), .SI(n33), .SE(reg_in[31]), .CK(clk), .Q(
        reg_out[31]) );
  SDFF_X1 reg_out_reg_30_ ( .D(1'b0), .SI(n33), .SE(reg_in[30]), .CK(clk), .Q(
        reg_out[30]) );
  SDFF_X1 reg_out_reg_29_ ( .D(1'b0), .SI(n33), .SE(reg_in[29]), .CK(clk), .Q(
        reg_out[29]) );
  SDFF_X1 reg_out_reg_28_ ( .D(1'b0), .SI(n33), .SE(reg_in[28]), .CK(clk), .Q(
        reg_out[28]) );
  SDFF_X1 reg_out_reg_27_ ( .D(1'b0), .SI(n33), .SE(reg_in[27]), .CK(clk), .Q(
        reg_out[27]) );
  SDFF_X1 reg_out_reg_26_ ( .D(1'b0), .SI(n33), .SE(reg_in[26]), .CK(clk), .Q(
        reg_out[26]) );
  SDFF_X1 reg_out_reg_25_ ( .D(1'b0), .SI(n33), .SE(reg_in[25]), .CK(clk), .Q(
        reg_out[25]) );
  SDFF_X1 reg_out_reg_24_ ( .D(1'b0), .SI(n33), .SE(reg_in[24]), .CK(clk), .Q(
        reg_out[24]) );
  SDFF_X1 reg_out_reg_23_ ( .D(1'b0), .SI(n33), .SE(reg_in[23]), .CK(clk), .Q(
        reg_out[23]) );
  SDFF_X1 reg_out_reg_22_ ( .D(1'b0), .SI(n33), .SE(reg_in[22]), .CK(clk), .Q(
        reg_out[22]) );
  SDFF_X1 reg_out_reg_21_ ( .D(1'b0), .SI(n33), .SE(reg_in[21]), .CK(clk), .Q(
        reg_out[21]) );
  SDFF_X1 reg_out_reg_20_ ( .D(1'b0), .SI(n34), .SE(reg_in[20]), .CK(clk), .Q(
        reg_out[20]) );
  SDFF_X1 reg_out_reg_19_ ( .D(1'b0), .SI(n34), .SE(reg_in[19]), .CK(clk), .Q(
        reg_out[19]) );
  SDFF_X1 reg_out_reg_18_ ( .D(1'b0), .SI(n34), .SE(reg_in[18]), .CK(clk), .Q(
        reg_out[18]) );
  SDFF_X1 reg_out_reg_17_ ( .D(1'b0), .SI(n34), .SE(reg_in[17]), .CK(clk), .Q(
        reg_out[17]) );
  SDFF_X1 reg_out_reg_16_ ( .D(1'b0), .SI(n34), .SE(reg_in[16]), .CK(clk), .Q(
        reg_out[16]) );
  SDFF_X1 reg_out_reg_15_ ( .D(1'b0), .SI(n34), .SE(reg_in[15]), .CK(clk), .Q(
        reg_out[15]) );
  SDFF_X1 reg_out_reg_14_ ( .D(1'b0), .SI(n34), .SE(reg_in[14]), .CK(clk), .Q(
        reg_out[14]) );
  SDFF_X1 reg_out_reg_13_ ( .D(1'b0), .SI(n34), .SE(reg_in[13]), .CK(clk), .Q(
        reg_out[13]) );
  SDFF_X1 reg_out_reg_12_ ( .D(1'b0), .SI(n34), .SE(reg_in[12]), .CK(clk), .Q(
        reg_out[12]) );
  SDFF_X1 reg_out_reg_11_ ( .D(1'b0), .SI(n34), .SE(reg_in[11]), .CK(clk), .Q(
        reg_out[11]) );
  SDFF_X1 reg_out_reg_10_ ( .D(1'b0), .SI(n34), .SE(reg_in[10]), .CK(clk), .Q(
        reg_out[10]) );
  SDFF_X1 reg_out_reg_9_ ( .D(1'b0), .SI(n35), .SE(reg_in[9]), .CK(clk), .Q(
        reg_out[9]) );
  SDFF_X1 reg_out_reg_8_ ( .D(1'b0), .SI(n35), .SE(reg_in[8]), .CK(clk), .Q(
        reg_out[8]) );
  SDFF_X1 reg_out_reg_7_ ( .D(1'b0), .SI(n35), .SE(reg_in[7]), .CK(clk), .Q(
        reg_out[7]) );
  SDFF_X1 reg_out_reg_6_ ( .D(1'b0), .SI(n35), .SE(reg_in[6]), .CK(clk), .Q(
        reg_out[6]) );
  SDFF_X1 reg_out_reg_5_ ( .D(1'b0), .SI(n35), .SE(reg_in[5]), .CK(clk), .Q(
        reg_out[5]) );
  SDFF_X1 reg_out_reg_4_ ( .D(1'b0), .SI(n35), .SE(reg_in[4]), .CK(clk), .Q(
        reg_out[4]) );
  SDFF_X1 reg_out_reg_3_ ( .D(1'b0), .SI(n35), .SE(reg_in[3]), .CK(clk), .Q(
        reg_out[3]) );
  SDFF_X1 reg_out_reg_2_ ( .D(1'b0), .SI(n35), .SE(reg_in[2]), .CK(clk), .Q(
        reg_out[2]) );
  SDFF_X1 reg_out_reg_1_ ( .D(1'b0), .SI(n35), .SE(reg_in[1]), .CK(clk), .Q(
        reg_out[1]) );
  SDFF_X1 reg_out_reg_0_ ( .D(1'b0), .SI(n35), .SE(reg_in[0]), .CK(clk), .Q(
        reg_out[0]) );
  BUF_X1 U35 ( .A(n36), .Z(n34) );
  BUF_X1 U36 ( .A(n36), .Z(n33) );
  BUF_X1 U37 ( .A(n36), .Z(n35) );
  INV_X1 U38 ( .A(reset), .ZN(n36) );
endmodule


module carryLookAheadAdder_0 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32;

  XOR2_X1 U66 ( .A(n24), .B(n35), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n36), .B(n25), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n26), .B(n37), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n38), .B(n27), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n28), .B(n39), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n40), .B(n29), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n41), .B(n42), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n43), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n30), .B(n44), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n45), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n46), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n47), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n48), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n49), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n50), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n51), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n52), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n53), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n54), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n55), .B(n31), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n56), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n57), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n58), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n59), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n60), .B(n17), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n18), .B(n61), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n62), .B(n19), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n20), .B(n63), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n64), .B(n21), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n22), .B(n65), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n66), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n32), .B(b[31]), .Z(n41) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n43) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n45) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n46) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n47) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n48) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n49) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n50) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n51) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n52) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n53) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n54) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n56) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n57) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n58) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n59) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n60) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n61) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n62) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n63) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n64) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n65) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n33) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n35) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n36) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n37) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n38) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n39) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n40) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n44) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n55) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n66) );
  INV_X1 U1 ( .A(n89), .ZN(n25) );
  AOI22_X1 U2 ( .A1(b[10]), .A2(a[10]), .B1(n22), .B2(n65), .ZN(n86) );
  INV_X1 U3 ( .A(n84), .ZN(n19) );
  AOI22_X1 U4 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n43), .ZN(n42) );
  INV_X1 U5 ( .A(n94), .ZN(n30) );
  OAI22_X1 U6 ( .A1(n1), .A2(n32), .B1(n42), .B2(n41), .ZN(cout) );
  INV_X1 U7 ( .A(b[31]), .ZN(n1) );
  INV_X1 U8 ( .A(n95), .ZN(n31) );
  AOI22_X1 U9 ( .A1(b[0]), .A2(a[0]), .B1(n66), .B2(cin), .ZN(n95) );
  INV_X1 U10 ( .A(a[31]), .ZN(n32) );
  AOI22_X1 U11 ( .A1(b[6]), .A2(a[6]), .B1(n26), .B2(n37), .ZN(n89) );
  AOI22_X1 U12 ( .A1(b[2]), .A2(a[2]), .B1(n30), .B2(n44), .ZN(n93) );
  INV_X1 U13 ( .A(n91), .ZN(n27) );
  AOI22_X1 U14 ( .A1(b[8]), .A2(a[8]), .B1(n24), .B2(n35), .ZN(n34) );
  INV_X1 U15 ( .A(n70), .ZN(n5) );
  INV_X1 U16 ( .A(n76), .ZN(n11) );
  AOI22_X1 U17 ( .A1(b[14]), .A2(a[14]), .B1(n18), .B2(n61), .ZN(n82) );
  AOI22_X1 U18 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n54), .ZN(n76) );
  AOI22_X1 U19 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n48), .ZN(n70) );
  AOI22_X1 U20 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n47), .ZN(n69) );
  AOI22_X1 U21 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n53), .ZN(n75) );
  AOI22_X1 U22 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n57), .ZN(n78) );
  AOI22_X1 U23 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n50), .ZN(n72) );
  AOI22_X1 U24 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n56), .ZN(n77) );
  AOI22_X1 U25 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n51), .ZN(n73) );
  AOI22_X1 U26 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n59), .ZN(n80) );
  AOI22_X1 U27 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n58), .ZN(n79) );
  AOI22_X1 U28 ( .A1(b[12]), .A2(a[12]), .B1(n20), .B2(n63), .ZN(n84) );
  AOI22_X1 U29 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n46), .ZN(n68) );
  INV_X1 U30 ( .A(n67), .ZN(n2) );
  AOI22_X1 U31 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n45), .ZN(n67) );
  AOI22_X1 U32 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n52), .ZN(n74) );
  INV_X1 U33 ( .A(n77), .ZN(n12) );
  INV_X1 U34 ( .A(n85), .ZN(n20) );
  INV_X1 U35 ( .A(n88), .ZN(n24) );
  AOI22_X1 U36 ( .A1(b[4]), .A2(a[4]), .B1(n28), .B2(n39), .ZN(n91) );
  INV_X1 U37 ( .A(n71), .ZN(n6) );
  AOI22_X1 U38 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n49), .ZN(n71) );
  INV_X1 U39 ( .A(n72), .ZN(n7) );
  AOI22_X1 U40 ( .A1(b[9]), .A2(a[9]), .B1(n23), .B2(n33), .ZN(n87) );
  AOI22_X1 U41 ( .A1(b[15]), .A2(a[15]), .B1(n17), .B2(n60), .ZN(n81) );
  AOI22_X1 U42 ( .A1(b[11]), .A2(a[11]), .B1(n21), .B2(n64), .ZN(n85) );
  INV_X1 U43 ( .A(n90), .ZN(n26) );
  INV_X1 U44 ( .A(n92), .ZN(n28) );
  AOI22_X1 U45 ( .A1(b[3]), .A2(a[3]), .B1(n29), .B2(n40), .ZN(n92) );
  AOI22_X1 U46 ( .A1(b[13]), .A2(a[13]), .B1(n19), .B2(n62), .ZN(n83) );
  AOI22_X1 U47 ( .A1(b[7]), .A2(a[7]), .B1(n25), .B2(n36), .ZN(n88) );
  INV_X1 U48 ( .A(n74), .ZN(n9) );
  INV_X1 U49 ( .A(n75), .ZN(n10) );
  INV_X1 U50 ( .A(n80), .ZN(n15) );
  INV_X1 U51 ( .A(n81), .ZN(n16) );
  INV_X1 U52 ( .A(n82), .ZN(n17) );
  INV_X1 U53 ( .A(n86), .ZN(n21) );
  AOI22_X1 U54 ( .A1(b[5]), .A2(a[5]), .B1(n27), .B2(n38), .ZN(n90) );
  INV_X1 U55 ( .A(n68), .ZN(n3) );
  INV_X1 U56 ( .A(n69), .ZN(n4) );
  INV_X1 U57 ( .A(n73), .ZN(n8) );
  INV_X1 U58 ( .A(n78), .ZN(n13) );
  INV_X1 U59 ( .A(n79), .ZN(n14) );
  INV_X1 U60 ( .A(n83), .ZN(n18) );
  INV_X1 U61 ( .A(n93), .ZN(n29) );
  INV_X1 U62 ( .A(n87), .ZN(n22) );
  XNOR2_X1 U63 ( .A(n33), .B(n34), .ZN(result[9]) );
  INV_X1 U64 ( .A(n34), .ZN(n23) );
  AOI22_X1 U65 ( .A1(b[1]), .A2(a[1]), .B1(n31), .B2(n55), .ZN(n94) );
endmodule


module carryLookAheadAdder_30 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n3), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n4), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n5), .B(n145), .Z(result[28]) );
  XOR2_X1 U78 ( .A(n7), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n8), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n9), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n10), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n11), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n12), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n13), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n14), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n15), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n16), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n17), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n2), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  INV_X1 U1 ( .A(n110), .ZN(n17) );
  INV_X1 U2 ( .A(n108), .ZN(n19) );
  INV_X1 U3 ( .A(n104), .ZN(n23) );
  AOI22_X1 U4 ( .A1(b[30]), .A2(a[30]), .B1(n3), .B2(n148), .ZN(n149) );
  INV_X1 U5 ( .A(n99), .ZN(n29) );
  OAI22_X1 U6 ( .A1(n1), .A2(n2), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U7 ( .A(b[31]), .ZN(n1) );
  INV_X1 U8 ( .A(a[31]), .ZN(n2) );
  INV_X1 U9 ( .A(n97), .ZN(n31) );
  INV_X1 U10 ( .A(n96), .ZN(n32) );
  AOI22_X1 U11 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U12 ( .A(n118), .ZN(n9) );
  INV_X1 U13 ( .A(n116), .ZN(n11) );
  INV_X1 U14 ( .A(n109), .ZN(n18) );
  INV_X1 U15 ( .A(n103), .ZN(n25) );
  XNOR2_X1 U16 ( .A(n144), .B(n121), .ZN(result[27]) );
  INV_X1 U17 ( .A(n122), .ZN(n5) );
  INV_X1 U18 ( .A(n124), .ZN(n3) );
  AOI22_X1 U19 ( .A1(b[29]), .A2(a[29]), .B1(n4), .B2(n146), .ZN(n124) );
  AOI22_X1 U20 ( .A1(b[25]), .A2(a[25]), .B1(n8), .B2(n142), .ZN(n120) );
  INV_X1 U21 ( .A(n106), .ZN(n21) );
  INV_X1 U22 ( .A(n100), .ZN(n28) );
  INV_X1 U23 ( .A(n101), .ZN(n27) );
  INV_X1 U24 ( .A(n112), .ZN(n15) );
  AOI22_X1 U25 ( .A1(b[24]), .A2(a[24]), .B1(n9), .B2(n141), .ZN(n119) );
  AOI22_X1 U26 ( .A1(b[27]), .A2(a[27]), .B1(n6), .B2(n144), .ZN(n122) );
  AOI22_X1 U27 ( .A1(b[21]), .A2(a[21]), .B1(n12), .B2(n138), .ZN(n116) );
  AOI22_X1 U28 ( .A1(b[23]), .A2(a[23]), .B1(n10), .B2(n140), .ZN(n118) );
  AOI22_X1 U29 ( .A1(b[26]), .A2(a[26]), .B1(n7), .B2(n143), .ZN(n121) );
  AOI22_X1 U30 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U31 ( .A1(b[28]), .A2(a[28]), .B1(n5), .B2(n145), .ZN(n123) );
  AOI22_X1 U32 ( .A1(b[22]), .A2(a[22]), .B1(n11), .B2(n139), .ZN(n117) );
  AOI22_X1 U33 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  AOI22_X1 U34 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
  INV_X1 U35 ( .A(n120), .ZN(n7) );
  AOI22_X1 U36 ( .A1(b[20]), .A2(a[20]), .B1(n13), .B2(n137), .ZN(n115) );
  AOI22_X1 U37 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U38 ( .A1(b[19]), .A2(a[19]), .B1(n14), .B2(n135), .ZN(n114) );
  AOI22_X1 U39 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  INV_X1 U40 ( .A(n98), .ZN(n30) );
  AOI22_X1 U41 ( .A1(b[17]), .A2(a[17]), .B1(n16), .B2(n133), .ZN(n112) );
  INV_X1 U42 ( .A(n123), .ZN(n4) );
  INV_X1 U43 ( .A(n121), .ZN(n6) );
  INV_X1 U44 ( .A(n119), .ZN(n8) );
  INV_X1 U45 ( .A(n114), .ZN(n13) );
  AOI22_X1 U46 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  AOI22_X1 U47 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  AOI22_X1 U48 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  AOI22_X1 U49 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U50 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  AOI22_X1 U51 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  AOI22_X1 U52 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U53 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U54 ( .A1(b[18]), .A2(a[18]), .B1(n15), .B2(n134), .ZN(n113) );
  AOI22_X1 U55 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  INV_X1 U56 ( .A(n117), .ZN(n10) );
  INV_X1 U57 ( .A(n115), .ZN(n12) );
  INV_X1 U58 ( .A(n113), .ZN(n14) );
  INV_X1 U59 ( .A(n111), .ZN(n16) );
  INV_X1 U60 ( .A(n107), .ZN(n20) );
  INV_X1 U61 ( .A(n105), .ZN(n22) );
  XNOR2_X1 U62 ( .A(n158), .B(n157), .ZN(result[9]) );
  INV_X1 U63 ( .A(n157), .ZN(n24) );
  INV_X1 U64 ( .A(n102), .ZN(n26) );
  AOI22_X1 U65 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U77 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
endmodule


module carryLookAheadAdder_29 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n3), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n4), .Z(result[29]) );
  XOR2_X1 U77 ( .A(n144), .B(n6), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n7), .B(n143), .Z(result[26]) );
  XOR2_X1 U80 ( .A(n9), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n10), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n11), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n12), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n13), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n14), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n15), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n16), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n17), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n2), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  INV_X1 U1 ( .A(n106), .ZN(n21) );
  INV_X1 U2 ( .A(n108), .ZN(n19) );
  INV_X1 U3 ( .A(b[31]), .ZN(n1) );
  INV_X1 U4 ( .A(n98), .ZN(n30) );
  INV_X1 U5 ( .A(a[31]), .ZN(n2) );
  INV_X1 U6 ( .A(n97), .ZN(n31) );
  INV_X1 U7 ( .A(n96), .ZN(n32) );
  AOI22_X1 U8 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U9 ( .A(n116), .ZN(n11) );
  OAI22_X1 U10 ( .A1(n1), .A2(n2), .B1(n149), .B2(n150), .ZN(cout) );
  AOI22_X1 U11 ( .A1(b[17]), .A2(a[17]), .B1(n16), .B2(n133), .ZN(n112) );
  INV_X1 U12 ( .A(n124), .ZN(n3) );
  AOI22_X1 U13 ( .A1(b[30]), .A2(a[30]), .B1(n3), .B2(n148), .ZN(n149) );
  AOI22_X1 U14 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  XNOR2_X1 U15 ( .A(n142), .B(n119), .ZN(result[25]) );
  XNOR2_X1 U16 ( .A(n122), .B(n145), .ZN(result[28]) );
  INV_X1 U17 ( .A(n123), .ZN(n4) );
  INV_X1 U18 ( .A(n120), .ZN(n7) );
  INV_X1 U19 ( .A(n118), .ZN(n9) );
  AOI22_X1 U20 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  AOI22_X1 U21 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  AOI22_X1 U22 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  INV_X1 U23 ( .A(n113), .ZN(n14) );
  AOI22_X1 U24 ( .A1(b[18]), .A2(a[18]), .B1(n15), .B2(n134), .ZN(n113) );
  INV_X1 U25 ( .A(n110), .ZN(n17) );
  AOI22_X1 U26 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U27 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  AOI22_X1 U28 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U29 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
  AOI22_X1 U30 ( .A1(b[22]), .A2(a[22]), .B1(n11), .B2(n139), .ZN(n117) );
  AOI22_X1 U31 ( .A1(b[26]), .A2(a[26]), .B1(n7), .B2(n143), .ZN(n121) );
  AOI22_X1 U32 ( .A1(b[29]), .A2(a[29]), .B1(n4), .B2(n146), .ZN(n124) );
  AOI22_X1 U33 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U34 ( .A1(b[20]), .A2(a[20]), .B1(n13), .B2(n137), .ZN(n115) );
  AOI22_X1 U35 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U36 ( .A1(b[28]), .A2(a[28]), .B1(n5), .B2(n145), .ZN(n123) );
  INV_X1 U37 ( .A(n119), .ZN(n8) );
  AOI22_X1 U38 ( .A1(b[24]), .A2(a[24]), .B1(n9), .B2(n141), .ZN(n119) );
  AOI22_X1 U39 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U40 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  INV_X1 U41 ( .A(n114), .ZN(n13) );
  INV_X1 U42 ( .A(n105), .ZN(n22) );
  INV_X1 U43 ( .A(n104), .ZN(n23) );
  INV_X1 U44 ( .A(n101), .ZN(n27) );
  AOI22_X1 U45 ( .A1(b[19]), .A2(a[19]), .B1(n14), .B2(n135), .ZN(n114) );
  AOI22_X1 U46 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  AOI22_X1 U47 ( .A1(b[21]), .A2(a[21]), .B1(n12), .B2(n138), .ZN(n116) );
  INV_X1 U48 ( .A(n115), .ZN(n12) );
  AOI22_X1 U49 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  INV_X1 U50 ( .A(n109), .ZN(n18) );
  INV_X1 U51 ( .A(n100), .ZN(n28) );
  AOI22_X1 U52 ( .A1(b[25]), .A2(a[25]), .B1(n8), .B2(n142), .ZN(n120) );
  INV_X1 U53 ( .A(n99), .ZN(n29) );
  AOI22_X1 U54 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U55 ( .A1(b[27]), .A2(a[27]), .B1(n6), .B2(n144), .ZN(n122) );
  INV_X1 U56 ( .A(n122), .ZN(n5) );
  INV_X1 U57 ( .A(n121), .ZN(n6) );
  AOI22_X1 U58 ( .A1(b[23]), .A2(a[23]), .B1(n10), .B2(n140), .ZN(n118) );
  INV_X1 U59 ( .A(n117), .ZN(n10) );
  INV_X1 U60 ( .A(n112), .ZN(n15) );
  INV_X1 U61 ( .A(n111), .ZN(n16) );
  INV_X1 U62 ( .A(n107), .ZN(n20) );
  XNOR2_X1 U63 ( .A(n158), .B(n157), .ZN(result[9]) );
  INV_X1 U64 ( .A(n157), .ZN(n24) );
  INV_X1 U65 ( .A(n103), .ZN(n25) );
  INV_X1 U76 ( .A(n102), .ZN(n26) );
  AOI22_X1 U79 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
endmodule


module carryLookAheadAdder_28 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n3), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n4), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n5), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n6), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n7), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n8), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n9), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n10), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n11), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n12), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n13), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n14), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n15), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n16), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n17), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n2), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  INV_X1 U1 ( .A(n110), .ZN(n17) );
  INV_X1 U2 ( .A(n104), .ZN(n23) );
  INV_X1 U3 ( .A(b[31]), .ZN(n1) );
  INV_X1 U4 ( .A(n102), .ZN(n26) );
  INV_X1 U5 ( .A(a[31]), .ZN(n2) );
  INV_X1 U6 ( .A(n99), .ZN(n29) );
  INV_X1 U7 ( .A(n96), .ZN(n32) );
  AOI22_X1 U8 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  AOI22_X1 U9 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  INV_X1 U10 ( .A(n108), .ZN(n19) );
  INV_X1 U11 ( .A(n122), .ZN(n5) );
  AOI22_X1 U12 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  OAI22_X1 U13 ( .A1(n1), .A2(n2), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U14 ( .A(n124), .ZN(n3) );
  AOI22_X1 U15 ( .A1(b[30]), .A2(a[30]), .B1(n3), .B2(n148), .ZN(n149) );
  INV_X1 U16 ( .A(n119), .ZN(n8) );
  INV_X1 U17 ( .A(n123), .ZN(n4) );
  AOI22_X1 U18 ( .A1(b[27]), .A2(a[27]), .B1(n6), .B2(n144), .ZN(n122) );
  AOI22_X1 U19 ( .A1(b[28]), .A2(a[28]), .B1(n5), .B2(n145), .ZN(n123) );
  XNOR2_X1 U20 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U21 ( .A1(b[24]), .A2(a[24]), .B1(n9), .B2(n141), .ZN(n119) );
  INV_X1 U22 ( .A(n118), .ZN(n9) );
  AOI22_X1 U23 ( .A1(b[23]), .A2(a[23]), .B1(n10), .B2(n140), .ZN(n118) );
  AOI22_X1 U24 ( .A1(b[22]), .A2(a[22]), .B1(n11), .B2(n139), .ZN(n117) );
  AOI22_X1 U25 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  INV_X1 U26 ( .A(n116), .ZN(n11) );
  INV_X1 U27 ( .A(n114), .ZN(n13) );
  AOI22_X1 U28 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U29 ( .A1(b[26]), .A2(a[26]), .B1(n7), .B2(n143), .ZN(n121) );
  AOI22_X1 U30 ( .A1(b[20]), .A2(a[20]), .B1(n13), .B2(n137), .ZN(n115) );
  AOI22_X1 U31 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  AOI22_X1 U32 ( .A1(b[17]), .A2(a[17]), .B1(n16), .B2(n133), .ZN(n112) );
  INV_X1 U33 ( .A(n105), .ZN(n22) );
  AOI22_X1 U34 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U35 ( .A1(b[19]), .A2(a[19]), .B1(n14), .B2(n135), .ZN(n114) );
  AOI22_X1 U36 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  INV_X1 U37 ( .A(n101), .ZN(n27) );
  INV_X1 U38 ( .A(n100), .ZN(n28) );
  AOI22_X1 U39 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  AOI22_X1 U40 ( .A1(b[29]), .A2(a[29]), .B1(n4), .B2(n146), .ZN(n124) );
  AOI22_X1 U41 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  INV_X1 U42 ( .A(n121), .ZN(n6) );
  INV_X1 U43 ( .A(n120), .ZN(n7) );
  INV_X1 U44 ( .A(n117), .ZN(n10) );
  AOI22_X1 U45 ( .A1(b[21]), .A2(a[21]), .B1(n12), .B2(n138), .ZN(n116) );
  INV_X1 U46 ( .A(n115), .ZN(n12) );
  INV_X1 U47 ( .A(n111), .ZN(n16) );
  INV_X1 U48 ( .A(n109), .ZN(n18) );
  INV_X1 U49 ( .A(n107), .ZN(n20) );
  AOI22_X1 U50 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U51 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U52 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
  INV_X1 U53 ( .A(n98), .ZN(n30) );
  INV_X1 U54 ( .A(n157), .ZN(n24) );
  AOI22_X1 U55 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  INV_X1 U56 ( .A(n113), .ZN(n14) );
  AOI22_X1 U57 ( .A1(b[18]), .A2(a[18]), .B1(n15), .B2(n134), .ZN(n113) );
  INV_X1 U58 ( .A(n112), .ZN(n15) );
  AOI22_X1 U59 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  INV_X1 U60 ( .A(n106), .ZN(n21) );
  AOI22_X1 U61 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  INV_X1 U62 ( .A(n97), .ZN(n31) );
  INV_X1 U63 ( .A(n103), .ZN(n25) );
  AOI22_X1 U64 ( .A1(b[25]), .A2(a[25]), .B1(n8), .B2(n142), .ZN(n120) );
  AOI22_X1 U65 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
endmodule


module carryLookAheadAdder_27 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n3), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n4), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n5), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n6), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n7), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n8), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n9), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n10), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n11), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n12), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n13), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n14), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n15), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n16), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n17), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n2), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  XOR2_X1 U1 ( .A(a[26]), .B(b[26]), .Z(n143) );
  INV_X1 U2 ( .A(n108), .ZN(n19) );
  INV_X1 U3 ( .A(n157), .ZN(n24) );
  INV_X1 U4 ( .A(b[31]), .ZN(n1) );
  INV_X1 U5 ( .A(a[31]), .ZN(n2) );
  INV_X1 U6 ( .A(n122), .ZN(n5) );
  INV_X1 U7 ( .A(n98), .ZN(n30) );
  INV_X1 U8 ( .A(n97), .ZN(n31) );
  INV_X1 U9 ( .A(n96), .ZN(n32) );
  AOI22_X1 U10 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U11 ( .A(n111), .ZN(n16) );
  AOI22_X1 U12 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  INV_X1 U13 ( .A(n118), .ZN(n9) );
  AOI22_X1 U14 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  INV_X1 U15 ( .A(n102), .ZN(n26) );
  INV_X1 U16 ( .A(n112), .ZN(n15) );
  OAI22_X1 U17 ( .A1(n1), .A2(n2), .B1(n149), .B2(n150), .ZN(cout) );
  AOI22_X1 U18 ( .A1(b[30]), .A2(a[30]), .B1(n3), .B2(n148), .ZN(n149) );
  INV_X1 U19 ( .A(n117), .ZN(n10) );
  INV_X1 U20 ( .A(n124), .ZN(n3) );
  AOI22_X1 U21 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  INV_X1 U22 ( .A(n109), .ZN(n18) );
  AOI22_X1 U23 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U24 ( .A1(b[18]), .A2(a[18]), .B1(n15), .B2(n134), .ZN(n113) );
  INV_X1 U25 ( .A(n123), .ZN(n4) );
  INV_X1 U26 ( .A(n119), .ZN(n8) );
  INV_X1 U27 ( .A(n116), .ZN(n11) );
  INV_X1 U28 ( .A(n114), .ZN(n13) );
  AOI22_X1 U29 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  AOI22_X1 U30 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  AOI22_X1 U31 ( .A1(b[28]), .A2(a[28]), .B1(n5), .B2(n145), .ZN(n123) );
  AOI22_X1 U32 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U33 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U34 ( .A1(b[29]), .A2(a[29]), .B1(n4), .B2(n146), .ZN(n124) );
  AOI22_X1 U35 ( .A1(b[24]), .A2(a[24]), .B1(n9), .B2(n141), .ZN(n119) );
  XNOR2_X1 U36 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U37 ( .A1(b[22]), .A2(a[22]), .B1(n11), .B2(n139), .ZN(n117) );
  AOI22_X1 U38 ( .A1(b[17]), .A2(a[17]), .B1(n16), .B2(n133), .ZN(n112) );
  AOI22_X1 U39 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  AOI22_X1 U40 ( .A1(b[21]), .A2(a[21]), .B1(n12), .B2(n138), .ZN(n116) );
  INV_X1 U41 ( .A(n121), .ZN(n6) );
  AOI22_X1 U42 ( .A1(b[26]), .A2(a[26]), .B1(n7), .B2(n143), .ZN(n121) );
  INV_X1 U43 ( .A(n115), .ZN(n12) );
  AOI22_X1 U44 ( .A1(b[20]), .A2(a[20]), .B1(n13), .B2(n137), .ZN(n115) );
  AOI22_X1 U45 ( .A1(b[19]), .A2(a[19]), .B1(n14), .B2(n135), .ZN(n114) );
  INV_X1 U46 ( .A(n120), .ZN(n7) );
  INV_X1 U47 ( .A(n107), .ZN(n20) );
  AOI22_X1 U48 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  INV_X1 U49 ( .A(n105), .ZN(n22) );
  INV_X1 U50 ( .A(n100), .ZN(n28) );
  INV_X1 U51 ( .A(n99), .ZN(n29) );
  AOI22_X1 U52 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U53 ( .A1(b[23]), .A2(a[23]), .B1(n10), .B2(n140), .ZN(n118) );
  AOI22_X1 U54 ( .A1(b[25]), .A2(a[25]), .B1(n8), .B2(n142), .ZN(n120) );
  AOI22_X1 U55 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U56 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
  INV_X1 U57 ( .A(n110), .ZN(n17) );
  AOI22_X1 U58 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  INV_X1 U59 ( .A(n104), .ZN(n23) );
  AOI22_X1 U60 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  INV_X1 U61 ( .A(n106), .ZN(n21) );
  AOI22_X1 U62 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  INV_X1 U63 ( .A(n101), .ZN(n27) );
  INV_X1 U64 ( .A(n103), .ZN(n25) );
  INV_X1 U65 ( .A(n113), .ZN(n14) );
  AOI22_X1 U102 ( .A1(b[27]), .A2(a[27]), .B1(n6), .B2(n144), .ZN(n122) );
endmodule


module carryLookAheadAdder_26 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n3), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n4), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n5), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n6), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n7), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n8), .Z(result[25]) );
  XOR2_X1 U81 ( .A(n140), .B(n10), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n11), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n12), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n13), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n14), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n15), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n16), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n17), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n2), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  OAI22_X1 U1 ( .A1(n1), .A2(n2), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U2 ( .A(b[31]), .ZN(n1) );
  INV_X1 U3 ( .A(a[31]), .ZN(n2) );
  INV_X1 U4 ( .A(n121), .ZN(n6) );
  INV_X1 U5 ( .A(n100), .ZN(n28) );
  INV_X1 U6 ( .A(n106), .ZN(n21) );
  INV_X1 U7 ( .A(n97), .ZN(n31) );
  INV_X1 U8 ( .A(n96), .ZN(n32) );
  AOI22_X1 U9 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U10 ( .A(n108), .ZN(n19) );
  AOI22_X1 U11 ( .A1(b[30]), .A2(a[30]), .B1(n3), .B2(n148), .ZN(n149) );
  INV_X1 U12 ( .A(n105), .ZN(n22) );
  INV_X1 U13 ( .A(n99), .ZN(n29) );
  INV_X1 U14 ( .A(n114), .ZN(n13) );
  XNOR2_X1 U15 ( .A(n118), .B(n141), .ZN(result[24]) );
  INV_X1 U16 ( .A(n120), .ZN(n7) );
  INV_X1 U17 ( .A(n98), .ZN(n30) );
  INV_X1 U18 ( .A(n123), .ZN(n4) );
  INV_X1 U19 ( .A(n117), .ZN(n10) );
  INV_X1 U20 ( .A(n112), .ZN(n15) );
  AOI22_X1 U21 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  INV_X1 U22 ( .A(n115), .ZN(n12) );
  AOI22_X1 U23 ( .A1(b[25]), .A2(a[25]), .B1(n8), .B2(n142), .ZN(n120) );
  AOI22_X1 U24 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  INV_X1 U25 ( .A(n119), .ZN(n8) );
  AOI22_X1 U26 ( .A1(b[26]), .A2(a[26]), .B1(n7), .B2(n143), .ZN(n121) );
  AOI22_X1 U27 ( .A1(b[19]), .A2(a[19]), .B1(n14), .B2(n135), .ZN(n114) );
  AOI22_X1 U28 ( .A1(b[22]), .A2(a[22]), .B1(n11), .B2(n139), .ZN(n117) );
  AOI22_X1 U29 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  XNOR2_X1 U30 ( .A(n158), .B(n157), .ZN(result[9]) );
  INV_X1 U31 ( .A(n157), .ZN(n24) );
  AOI22_X1 U32 ( .A1(b[20]), .A2(a[20]), .B1(n13), .B2(n137), .ZN(n115) );
  INV_X1 U33 ( .A(n124), .ZN(n3) );
  AOI22_X1 U34 ( .A1(b[29]), .A2(a[29]), .B1(n4), .B2(n146), .ZN(n124) );
  AOI22_X1 U35 ( .A1(b[18]), .A2(a[18]), .B1(n15), .B2(n134), .ZN(n113) );
  AOI22_X1 U36 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U37 ( .A1(b[28]), .A2(a[28]), .B1(n5), .B2(n145), .ZN(n123) );
  AOI22_X1 U38 ( .A1(b[24]), .A2(a[24]), .B1(n9), .B2(n141), .ZN(n119) );
  INV_X1 U39 ( .A(n109), .ZN(n18) );
  INV_X1 U40 ( .A(n122), .ZN(n5) );
  INV_X1 U41 ( .A(n118), .ZN(n9) );
  INV_X1 U42 ( .A(n116), .ZN(n11) );
  INV_X1 U43 ( .A(n113), .ZN(n14) );
  AOI22_X1 U44 ( .A1(b[17]), .A2(a[17]), .B1(n16), .B2(n133), .ZN(n112) );
  AOI22_X1 U45 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  AOI22_X1 U46 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  INV_X1 U47 ( .A(n107), .ZN(n20) );
  AOI22_X1 U48 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U49 ( .A1(b[27]), .A2(a[27]), .B1(n6), .B2(n144), .ZN(n122) );
  AOI22_X1 U50 ( .A1(b[21]), .A2(a[21]), .B1(n12), .B2(n138), .ZN(n116) );
  AOI22_X1 U51 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U52 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U53 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U54 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  AOI22_X1 U55 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  INV_X1 U56 ( .A(n111), .ZN(n16) );
  AOI22_X1 U57 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
  INV_X1 U58 ( .A(n102), .ZN(n26) );
  AOI22_X1 U59 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  INV_X1 U60 ( .A(n110), .ZN(n17) );
  AOI22_X1 U61 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  INV_X1 U62 ( .A(n104), .ZN(n23) );
  INV_X1 U63 ( .A(n101), .ZN(n27) );
  AOI22_X1 U64 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  INV_X1 U65 ( .A(n103), .ZN(n25) );
  AOI22_X1 U80 ( .A1(b[23]), .A2(a[23]), .B1(n10), .B2(n140), .ZN(n118) );
endmodule


module carryLookAheadAdder_25 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159;

  XOR2_X1 U66 ( .A(n26), .B(n157), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n156), .B(n27), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n28), .B(n155), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n154), .B(n29), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n30), .B(n153), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n152), .B(n31), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n151), .B(n150), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n4), .B(n149), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n32), .B(n148), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n147), .B(n5), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n6), .B(n146), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n145), .B(n7), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n8), .B(n144), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n143), .B(n9), .Z(result[25]) );
  XOR2_X1 U81 ( .A(n141), .B(n11), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n12), .B(n140), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n139), .B(n13), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n14), .B(n138), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n137), .B(n96), .Z(result[1]) );
  XOR2_X1 U87 ( .A(n16), .B(n135), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n134), .B(n17), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n18), .B(n133), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n132), .B(n19), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n20), .B(n131), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n130), .B(n21), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n22), .B(n129), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n128), .B(n23), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n24), .B(n127), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n126), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n3), .B(b[31]), .Z(n151) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n149) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n147) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n146) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n145) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n144) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n143) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n142) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n139) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n138) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n136) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n135) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n134) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n133) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n132) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n131) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n130) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n129) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n128) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n127) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n159) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n157) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n156) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n155) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n154) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n153) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n152) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n148) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n137) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n126) );
  XOR2_X1 U1 ( .A(a[22]), .B(b[22]), .Z(n140) );
  INV_X1 U2 ( .A(b[23]), .ZN(n1) );
  INV_X1 U3 ( .A(n109), .ZN(n20) );
  INV_X1 U4 ( .A(a[31]), .ZN(n3) );
  INV_X1 U5 ( .A(b[31]), .ZN(n2) );
  INV_X1 U6 ( .A(n105), .ZN(n24) );
  INV_X1 U7 ( .A(n98), .ZN(n32) );
  INV_X1 U8 ( .A(n97), .ZN(n96) );
  AOI22_X1 U9 ( .A1(b[0]), .A2(a[0]), .B1(n126), .B2(cin), .ZN(n97) );
  INV_X1 U10 ( .A(n115), .ZN(n14) );
  INV_X1 U11 ( .A(n104), .ZN(n26) );
  INV_X1 U12 ( .A(n117), .ZN(n12) );
  XNOR2_X1 U13 ( .A(n119), .B(n142), .ZN(result[24]) );
  XNOR2_X1 U14 ( .A(n136), .B(n114), .ZN(result[19]) );
  INV_X1 U15 ( .A(n100), .ZN(n30) );
  XNOR2_X1 U16 ( .A(a[23]), .B(n1), .ZN(n141) );
  OAI22_X1 U17 ( .A1(n2), .A2(n3), .B1(n150), .B2(n151), .ZN(cout) );
  AOI22_X1 U18 ( .A1(b[30]), .A2(a[30]), .B1(n4), .B2(n149), .ZN(n150) );
  INV_X1 U19 ( .A(n122), .ZN(n7) );
  INV_X1 U20 ( .A(n119), .ZN(n10) );
  INV_X1 U21 ( .A(n113), .ZN(n16) );
  INV_X1 U22 ( .A(n102), .ZN(n28) );
  INV_X1 U23 ( .A(n125), .ZN(n4) );
  AOI22_X1 U24 ( .A1(b[23]), .A2(a[23]), .B1(n11), .B2(n141), .ZN(n119) );
  INV_X1 U25 ( .A(n124), .ZN(n5) );
  INV_X1 U26 ( .A(n118), .ZN(n11) );
  AOI22_X1 U27 ( .A1(b[6]), .A2(a[6]), .B1(n28), .B2(n155), .ZN(n103) );
  INV_X1 U28 ( .A(n112), .ZN(n17) );
  AOI22_X1 U29 ( .A1(b[5]), .A2(a[5]), .B1(n29), .B2(n154), .ZN(n102) );
  AOI22_X1 U30 ( .A1(b[4]), .A2(a[4]), .B1(n30), .B2(n153), .ZN(n101) );
  AOI22_X1 U31 ( .A1(b[8]), .A2(a[8]), .B1(n26), .B2(n157), .ZN(n158) );
  INV_X1 U32 ( .A(n123), .ZN(n6) );
  AOI22_X1 U33 ( .A1(b[18]), .A2(a[18]), .B1(n16), .B2(n135), .ZN(n114) );
  AOI22_X1 U34 ( .A1(b[10]), .A2(a[10]), .B1(n24), .B2(n127), .ZN(n106) );
  AOI22_X1 U35 ( .A1(b[22]), .A2(a[22]), .B1(n12), .B2(n140), .ZN(n118) );
  AOI22_X1 U36 ( .A1(b[2]), .A2(a[2]), .B1(n32), .B2(n148), .ZN(n99) );
  AOI22_X1 U37 ( .A1(b[21]), .A2(a[21]), .B1(n13), .B2(n139), .ZN(n117) );
  AOI22_X1 U38 ( .A1(b[11]), .A2(a[11]), .B1(n23), .B2(n128), .ZN(n107) );
  AOI22_X1 U39 ( .A1(b[29]), .A2(a[29]), .B1(n5), .B2(n147), .ZN(n125) );
  AOI22_X1 U40 ( .A1(b[14]), .A2(a[14]), .B1(n20), .B2(n131), .ZN(n110) );
  AOI22_X1 U41 ( .A1(b[20]), .A2(a[20]), .B1(n14), .B2(n138), .ZN(n116) );
  AOI22_X1 U42 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(n152), .ZN(n100) );
  AOI22_X1 U43 ( .A1(b[17]), .A2(a[17]), .B1(n17), .B2(n134), .ZN(n113) );
  AOI22_X1 U44 ( .A1(b[13]), .A2(a[13]), .B1(n21), .B2(n130), .ZN(n109) );
  AOI22_X1 U45 ( .A1(b[28]), .A2(a[28]), .B1(n6), .B2(n146), .ZN(n124) );
  AOI22_X1 U46 ( .A1(b[24]), .A2(a[24]), .B1(n10), .B2(n142), .ZN(n120) );
  INV_X1 U47 ( .A(n120), .ZN(n9) );
  INV_X1 U48 ( .A(n99), .ZN(n31) );
  AOI22_X1 U49 ( .A1(b[15]), .A2(a[15]), .B1(n19), .B2(n132), .ZN(n111) );
  AOI22_X1 U50 ( .A1(b[19]), .A2(a[19]), .B1(n15), .B2(n136), .ZN(n115) );
  AOI22_X1 U51 ( .A1(b[16]), .A2(a[16]), .B1(n18), .B2(n133), .ZN(n112) );
  INV_X1 U52 ( .A(n107), .ZN(n22) );
  INV_X1 U53 ( .A(n103), .ZN(n27) );
  AOI22_X1 U54 ( .A1(b[27]), .A2(a[27]), .B1(n7), .B2(n145), .ZN(n123) );
  AOI22_X1 U55 ( .A1(b[12]), .A2(a[12]), .B1(n22), .B2(n129), .ZN(n108) );
  AOI22_X1 U56 ( .A1(b[26]), .A2(a[26]), .B1(n8), .B2(n144), .ZN(n122) );
  INV_X1 U57 ( .A(n121), .ZN(n8) );
  INV_X1 U58 ( .A(n116), .ZN(n13) );
  INV_X1 U59 ( .A(n114), .ZN(n15) );
  INV_X1 U60 ( .A(n111), .ZN(n18) );
  AOI22_X1 U61 ( .A1(b[9]), .A2(a[9]), .B1(n25), .B2(n159), .ZN(n105) );
  AOI22_X1 U62 ( .A1(b[7]), .A2(a[7]), .B1(n27), .B2(n156), .ZN(n104) );
  INV_X1 U63 ( .A(n110), .ZN(n19) );
  INV_X1 U64 ( .A(n108), .ZN(n21) );
  INV_X1 U65 ( .A(n106), .ZN(n23) );
  XNOR2_X1 U80 ( .A(n159), .B(n158), .ZN(result[9]) );
  INV_X1 U86 ( .A(n158), .ZN(n25) );
  INV_X1 U105 ( .A(n101), .ZN(n29) );
  AOI22_X1 U106 ( .A1(b[1]), .A2(a[1]), .B1(n96), .B2(n137), .ZN(n98) );
  AOI22_X1 U129 ( .A1(b[25]), .A2(a[25]), .B1(n9), .B2(n143), .ZN(n121) );
endmodule


module carryLookAheadAdder_24 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n3), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n4), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n5), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n6), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n7), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n8), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n9), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n10), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n11), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n12), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n13), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n14), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n15), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n16), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n17), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n2), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  INV_X1 U1 ( .A(a[31]), .ZN(n2) );
  INV_X1 U2 ( .A(n100), .ZN(n28) );
  INV_X1 U3 ( .A(n103), .ZN(n25) );
  INV_X1 U4 ( .A(n106), .ZN(n21) );
  OAI22_X1 U5 ( .A1(n1), .A2(n2), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U6 ( .A(b[31]), .ZN(n1) );
  INV_X1 U7 ( .A(n99), .ZN(n29) );
  INV_X1 U8 ( .A(n96), .ZN(n32) );
  AOI22_X1 U9 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U10 ( .A(n114), .ZN(n13) );
  INV_X1 U11 ( .A(n104), .ZN(n23) );
  INV_X1 U12 ( .A(n113), .ZN(n14) );
  INV_X1 U13 ( .A(n98), .ZN(n30) );
  INV_X1 U14 ( .A(n120), .ZN(n7) );
  INV_X1 U15 ( .A(n122), .ZN(n5) );
  AOI22_X1 U16 ( .A1(b[20]), .A2(a[20]), .B1(n13), .B2(n137), .ZN(n115) );
  INV_X1 U17 ( .A(n97), .ZN(n31) );
  INV_X1 U18 ( .A(n101), .ZN(n27) );
  INV_X1 U19 ( .A(n110), .ZN(n17) );
  AOI22_X1 U20 ( .A1(b[21]), .A2(a[21]), .B1(n12), .B2(n138), .ZN(n116) );
  AOI22_X1 U21 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  INV_X1 U22 ( .A(n123), .ZN(n4) );
  AOI22_X1 U23 ( .A1(b[26]), .A2(a[26]), .B1(n7), .B2(n143), .ZN(n121) );
  INV_X1 U24 ( .A(n109), .ZN(n18) );
  INV_X1 U25 ( .A(n108), .ZN(n19) );
  AOI22_X1 U26 ( .A1(b[19]), .A2(a[19]), .B1(n14), .B2(n135), .ZN(n114) );
  AOI22_X1 U27 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  AOI22_X1 U28 ( .A1(b[30]), .A2(a[30]), .B1(n3), .B2(n148), .ZN(n149) );
  AOI22_X1 U29 ( .A1(b[28]), .A2(a[28]), .B1(n5), .B2(n145), .ZN(n123) );
  AOI22_X1 U30 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  AOI22_X1 U31 ( .A1(b[24]), .A2(a[24]), .B1(n9), .B2(n141), .ZN(n119) );
  INV_X1 U32 ( .A(n124), .ZN(n3) );
  INV_X1 U33 ( .A(n118), .ZN(n9) );
  INV_X1 U34 ( .A(n117), .ZN(n10) );
  AOI22_X1 U35 ( .A1(b[18]), .A2(a[18]), .B1(n15), .B2(n134), .ZN(n113) );
  INV_X1 U36 ( .A(n112), .ZN(n15) );
  INV_X1 U37 ( .A(n107), .ZN(n20) );
  AOI22_X1 U38 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U39 ( .A1(b[23]), .A2(a[23]), .B1(n10), .B2(n140), .ZN(n118) );
  INV_X1 U40 ( .A(n119), .ZN(n8) );
  AOI22_X1 U41 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U42 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U43 ( .A1(b[22]), .A2(a[22]), .B1(n11), .B2(n139), .ZN(n117) );
  AOI22_X1 U44 ( .A1(b[29]), .A2(a[29]), .B1(n4), .B2(n146), .ZN(n124) );
  AOI22_X1 U45 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  AOI22_X1 U46 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  AOI22_X1 U47 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U48 ( .A1(b[25]), .A2(a[25]), .B1(n8), .B2(n142), .ZN(n120) );
  AOI22_X1 U49 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  AOI22_X1 U50 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U51 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U52 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  AOI22_X1 U53 ( .A1(b[27]), .A2(a[27]), .B1(n6), .B2(n144), .ZN(n122) );
  INV_X1 U54 ( .A(n121), .ZN(n6) );
  INV_X1 U55 ( .A(n116), .ZN(n11) );
  INV_X1 U56 ( .A(n115), .ZN(n12) );
  AOI22_X1 U57 ( .A1(b[17]), .A2(a[17]), .B1(n16), .B2(n133), .ZN(n112) );
  INV_X1 U58 ( .A(n111), .ZN(n16) );
  INV_X1 U59 ( .A(n105), .ZN(n22) );
  XNOR2_X1 U60 ( .A(n158), .B(n157), .ZN(result[9]) );
  INV_X1 U61 ( .A(n157), .ZN(n24) );
  AOI22_X1 U62 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  INV_X1 U63 ( .A(n102), .ZN(n26) );
  AOI22_X1 U64 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U65 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
endmodule


module carryLookAheadAdder_23 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160;

  XOR2_X1 U66 ( .A(n27), .B(n158), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n157), .B(n28), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n29), .B(n156), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n155), .B(n30), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n31), .B(n154), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n153), .B(n32), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n152), .B(n151), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n5), .B(n150), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n96), .B(n149), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n148), .B(n6), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n7), .B(n147), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n146), .B(n8), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n9), .B(n145), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n144), .B(n10), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n11), .B(n143), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n142), .B(n12), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n13), .B(n141), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n140), .B(n14), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n15), .B(n139), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n138), .B(n97), .Z(result[1]) );
  XOR2_X1 U87 ( .A(n17), .B(n136), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n135), .B(n18), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n19), .B(n134), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n133), .B(n20), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n21), .B(n132), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n131), .B(n22), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n23), .B(n130), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n129), .B(n24), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n25), .B(n128), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n127), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n4), .B(b[31]), .Z(n152) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n150) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n148) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n147) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n146) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n145) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n144) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n143) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n142) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n140) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n137) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n135) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n134) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n133) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n132) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n131) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n130) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n129) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n128) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n160) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n158) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n157) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n156) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n155) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n154) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n153) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n149) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n138) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n127) );
  INV_X1 U1 ( .A(b[18]), .ZN(n1) );
  INV_X1 U2 ( .A(b[20]), .ZN(n2) );
  XOR2_X1 U3 ( .A(a[22]), .B(b[22]), .Z(n141) );
  INV_X1 U4 ( .A(b[31]), .ZN(n3) );
  INV_X1 U5 ( .A(n104), .ZN(n28) );
  INV_X1 U6 ( .A(a[31]), .ZN(n4) );
  INV_X1 U7 ( .A(n99), .ZN(n96) );
  INV_X1 U8 ( .A(n98), .ZN(n97) );
  AOI22_X1 U9 ( .A1(b[0]), .A2(a[0]), .B1(n127), .B2(cin), .ZN(n98) );
  INV_X1 U10 ( .A(n126), .ZN(n5) );
  AOI22_X1 U11 ( .A1(b[15]), .A2(a[15]), .B1(n20), .B2(n133), .ZN(n112) );
  XNOR2_X1 U12 ( .A(a[18]), .B(n1), .ZN(n136) );
  INV_X1 U13 ( .A(n112), .ZN(n19) );
  XNOR2_X1 U14 ( .A(a[20]), .B(n2), .ZN(n139) );
  XNOR2_X1 U15 ( .A(n137), .B(n115), .ZN(result[19]) );
  INV_X1 U16 ( .A(n114), .ZN(n17) );
  INV_X1 U17 ( .A(n108), .ZN(n23) );
  INV_X1 U18 ( .A(n103), .ZN(n29) );
  INV_X1 U19 ( .A(n124), .ZN(n7) );
  INV_X1 U20 ( .A(n121), .ZN(n10) );
  INV_X1 U21 ( .A(n120), .ZN(n11) );
  INV_X1 U22 ( .A(n105), .ZN(n27) );
  AOI22_X1 U23 ( .A1(b[24]), .A2(a[24]), .B1(n11), .B2(n143), .ZN(n121) );
  INV_X1 U24 ( .A(n110), .ZN(n21) );
  AOI22_X1 U25 ( .A1(b[12]), .A2(a[12]), .B1(n23), .B2(n130), .ZN(n109) );
  INV_X1 U26 ( .A(n107), .ZN(n24) );
  INV_X1 U27 ( .A(n101), .ZN(n31) );
  AOI22_X1 U28 ( .A1(b[2]), .A2(a[2]), .B1(n96), .B2(n149), .ZN(n100) );
  OAI22_X1 U29 ( .A1(n3), .A2(n4), .B1(n151), .B2(n152), .ZN(cout) );
  INV_X1 U30 ( .A(n123), .ZN(n8) );
  INV_X1 U31 ( .A(n119), .ZN(n12) );
  INV_X1 U32 ( .A(n117), .ZN(n14) );
  INV_X1 U33 ( .A(n113), .ZN(n18) );
  AOI22_X1 U34 ( .A1(b[11]), .A2(a[11]), .B1(n24), .B2(n129), .ZN(n108) );
  AOI22_X1 U35 ( .A1(b[23]), .A2(a[23]), .B1(n12), .B2(n142), .ZN(n120) );
  AOI22_X1 U36 ( .A1(b[13]), .A2(a[13]), .B1(n22), .B2(n131), .ZN(n110) );
  AOI22_X1 U37 ( .A1(b[16]), .A2(a[16]), .B1(n19), .B2(n134), .ZN(n113) );
  AOI22_X1 U38 ( .A1(b[8]), .A2(a[8]), .B1(n27), .B2(n158), .ZN(n159) );
  INV_X1 U39 ( .A(n102), .ZN(n30) );
  AOI22_X1 U40 ( .A1(b[1]), .A2(a[1]), .B1(n97), .B2(n138), .ZN(n99) );
  AOI22_X1 U41 ( .A1(b[28]), .A2(a[28]), .B1(n7), .B2(n147), .ZN(n125) );
  AOI22_X1 U42 ( .A1(b[14]), .A2(a[14]), .B1(n21), .B2(n132), .ZN(n111) );
  AOI22_X1 U43 ( .A1(b[18]), .A2(a[18]), .B1(n17), .B2(n136), .ZN(n115) );
  AOI22_X1 U44 ( .A1(b[4]), .A2(a[4]), .B1(n31), .B2(n154), .ZN(n102) );
  AOI22_X1 U45 ( .A1(b[30]), .A2(a[30]), .B1(n5), .B2(n150), .ZN(n151) );
  AOI22_X1 U46 ( .A1(b[27]), .A2(a[27]), .B1(n8), .B2(n146), .ZN(n124) );
  AOI22_X1 U47 ( .A1(b[26]), .A2(a[26]), .B1(n9), .B2(n145), .ZN(n123) );
  INV_X1 U48 ( .A(n122), .ZN(n9) );
  AOI22_X1 U49 ( .A1(b[20]), .A2(a[20]), .B1(n15), .B2(n139), .ZN(n117) );
  AOI22_X1 U50 ( .A1(b[10]), .A2(a[10]), .B1(n25), .B2(n128), .ZN(n107) );
  AOI22_X1 U51 ( .A1(b[5]), .A2(a[5]), .B1(n30), .B2(n155), .ZN(n103) );
  AOI22_X1 U52 ( .A1(b[3]), .A2(a[3]), .B1(n32), .B2(n153), .ZN(n101) );
  AOI22_X1 U53 ( .A1(b[22]), .A2(a[22]), .B1(n13), .B2(n141), .ZN(n119) );
  INV_X1 U54 ( .A(n125), .ZN(n6) );
  AOI22_X1 U55 ( .A1(b[17]), .A2(a[17]), .B1(n18), .B2(n135), .ZN(n114) );
  AOI22_X1 U56 ( .A1(b[25]), .A2(a[25]), .B1(n10), .B2(n144), .ZN(n122) );
  AOI22_X1 U57 ( .A1(b[6]), .A2(a[6]), .B1(n29), .B2(n156), .ZN(n104) );
  AOI22_X1 U58 ( .A1(b[7]), .A2(a[7]), .B1(n28), .B2(n157), .ZN(n105) );
  INV_X1 U59 ( .A(n118), .ZN(n13) );
  INV_X1 U60 ( .A(n116), .ZN(n15) );
  INV_X1 U61 ( .A(n115), .ZN(n16) );
  INV_X1 U62 ( .A(n111), .ZN(n20) );
  INV_X1 U63 ( .A(n109), .ZN(n22) );
  INV_X1 U64 ( .A(n106), .ZN(n25) );
  XNOR2_X1 U65 ( .A(n160), .B(n159), .ZN(result[9]) );
  INV_X1 U86 ( .A(n159), .ZN(n26) );
  AOI22_X1 U106 ( .A1(b[19]), .A2(a[19]), .B1(n16), .B2(n137), .ZN(n116) );
  INV_X1 U108 ( .A(n100), .ZN(n32) );
  AOI22_X1 U110 ( .A1(b[21]), .A2(a[21]), .B1(n14), .B2(n140), .ZN(n118) );
  AOI22_X1 U129 ( .A1(b[29]), .A2(a[29]), .B1(n6), .B2(n148), .ZN(n126) );
  AOI22_X1 U130 ( .A1(b[9]), .A2(a[9]), .B1(n26), .B2(n160), .ZN(n106) );
endmodule


module carryLookAheadAdder_22 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n3), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n4), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n5), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n6), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n7), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n8), .B(n142), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n9), .B(n141), .Z(result[24]) );
  XOR2_X1 U82 ( .A(n11), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n12), .B(n138), .Z(result[21]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n14), .B(n135), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n15), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n16), .Z(result[17]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n2), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  INV_X1 U1 ( .A(b[31]), .ZN(n1) );
  INV_X1 U2 ( .A(a[31]), .ZN(n2) );
  INV_X1 U3 ( .A(n101), .ZN(n27) );
  INV_X1 U4 ( .A(n99), .ZN(n29) );
  INV_X1 U5 ( .A(n97), .ZN(n31) );
  INV_X1 U6 ( .A(n96), .ZN(n32) );
  AOI22_X1 U7 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U8 ( .A(n104), .ZN(n23) );
  XNOR2_X1 U9 ( .A(n110), .B(n132), .ZN(result[16]) );
  INV_X1 U10 ( .A(n123), .ZN(n4) );
  XNOR2_X1 U11 ( .A(n140), .B(n117), .ZN(result[23]) );
  XNOR2_X1 U12 ( .A(n109), .B(n131), .ZN(result[15]) );
  XNOR2_X1 U13 ( .A(n114), .B(n137), .ZN(result[20]) );
  INV_X1 U14 ( .A(n116), .ZN(n11) );
  AOI22_X1 U15 ( .A1(b[28]), .A2(a[28]), .B1(n5), .B2(n145), .ZN(n123) );
  INV_X1 U16 ( .A(n103), .ZN(n25) );
  OAI22_X1 U17 ( .A1(n1), .A2(n2), .B1(n149), .B2(n150), .ZN(cout) );
  AOI22_X1 U18 ( .A1(b[30]), .A2(a[30]), .B1(n3), .B2(n148), .ZN(n149) );
  AOI22_X1 U19 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  INV_X1 U20 ( .A(n124), .ZN(n3) );
  INV_X1 U21 ( .A(n106), .ZN(n21) );
  INV_X1 U22 ( .A(n108), .ZN(n19) );
  AOI22_X1 U23 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  INV_X1 U24 ( .A(n122), .ZN(n5) );
  INV_X1 U25 ( .A(n118), .ZN(n9) );
  INV_X1 U26 ( .A(n115), .ZN(n12) );
  INV_X1 U27 ( .A(n112), .ZN(n15) );
  INV_X1 U28 ( .A(n110), .ZN(n17) );
  AOI22_X1 U29 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U30 ( .A1(b[21]), .A2(a[21]), .B1(n12), .B2(n138), .ZN(n116) );
  AOI22_X1 U31 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  AOI22_X1 U32 ( .A1(b[23]), .A2(a[23]), .B1(n10), .B2(n140), .ZN(n118) );
  AOI22_X1 U33 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  AOI22_X1 U34 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  AOI22_X1 U35 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  INV_X1 U36 ( .A(n102), .ZN(n26) );
  AOI22_X1 U37 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U38 ( .A1(b[20]), .A2(a[20]), .B1(n13), .B2(n137), .ZN(n115) );
  AOI22_X1 U39 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  INV_X1 U40 ( .A(n120), .ZN(n7) );
  INV_X1 U41 ( .A(n113), .ZN(n14) );
  AOI22_X1 U42 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
  AOI22_X1 U43 ( .A1(b[22]), .A2(a[22]), .B1(n11), .B2(n139), .ZN(n117) );
  AOI22_X1 U44 ( .A1(b[18]), .A2(a[18]), .B1(n15), .B2(n134), .ZN(n113) );
  AOI22_X1 U45 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  AOI22_X1 U46 ( .A1(b[29]), .A2(a[29]), .B1(n4), .B2(n146), .ZN(n124) );
  AOI22_X1 U47 ( .A1(b[26]), .A2(a[26]), .B1(n7), .B2(n143), .ZN(n121) );
  AOI22_X1 U48 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U49 ( .A1(b[27]), .A2(a[27]), .B1(n6), .B2(n144), .ZN(n122) );
  AOI22_X1 U50 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  AOI22_X1 U51 ( .A1(b[25]), .A2(a[25]), .B1(n8), .B2(n142), .ZN(n120) );
  AOI22_X1 U52 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U53 ( .A1(b[17]), .A2(a[17]), .B1(n16), .B2(n133), .ZN(n112) );
  AOI22_X1 U54 ( .A1(b[24]), .A2(a[24]), .B1(n9), .B2(n141), .ZN(n119) );
  INV_X1 U55 ( .A(n98), .ZN(n30) );
  INV_X1 U56 ( .A(n121), .ZN(n6) );
  INV_X1 U57 ( .A(n119), .ZN(n8) );
  INV_X1 U58 ( .A(n117), .ZN(n10) );
  INV_X1 U59 ( .A(n114), .ZN(n13) );
  INV_X1 U60 ( .A(n111), .ZN(n16) );
  INV_X1 U61 ( .A(n109), .ZN(n18) );
  INV_X1 U62 ( .A(n107), .ZN(n20) );
  INV_X1 U63 ( .A(n105), .ZN(n22) );
  XNOR2_X1 U64 ( .A(n158), .B(n157), .ZN(result[9]) );
  INV_X1 U65 ( .A(n157), .ZN(n24) );
  INV_X1 U81 ( .A(n100), .ZN(n28) );
  AOI22_X1 U84 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U89 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U90 ( .A1(b[19]), .A2(a[19]), .B1(n14), .B2(n135), .ZN(n114) );
endmodule


module carryLookAheadAdder_21 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159;

  XOR2_X1 U66 ( .A(n26), .B(n157), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n156), .B(n27), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n28), .B(n155), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n154), .B(n29), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n30), .B(n153), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n152), .B(n31), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n151), .B(n150), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n3), .B(n149), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n32), .B(n148), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n147), .B(n4), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n5), .B(n146), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n145), .B(n6), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n7), .B(n144), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n143), .B(n8), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n9), .B(n142), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n141), .B(n10), .Z(result[23]) );
  XOR2_X1 U83 ( .A(n139), .B(n13), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n14), .B(n138), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n137), .B(n96), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n136), .B(n15), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n16), .B(n135), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n134), .B(n17), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n18), .B(n133), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n132), .B(n19), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n20), .B(n131), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n130), .B(n21), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n22), .B(n129), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n128), .B(n23), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n24), .B(n127), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n126), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n2), .B(b[31]), .Z(n151) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n149) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n147) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n146) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n145) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n144) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n143) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n142) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n141) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n140) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n139) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n138) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n136) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n135) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n134) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n132) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n131) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n130) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n129) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n128) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n127) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n159) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n157) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n156) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n155) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n154) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n153) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n152) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n148) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n137) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n126) );
  INV_X1 U1 ( .A(b[16]), .ZN(n1) );
  INV_X1 U2 ( .A(b[31]), .ZN(n11) );
  INV_X1 U3 ( .A(a[31]), .ZN(n2) );
  INV_X1 U4 ( .A(n100), .ZN(n30) );
  INV_X1 U5 ( .A(n98), .ZN(n32) );
  INV_X1 U6 ( .A(n97), .ZN(n96) );
  AOI22_X1 U7 ( .A1(b[0]), .A2(a[0]), .B1(n126), .B2(cin), .ZN(n97) );
  XNOR2_X1 U8 ( .A(a[16]), .B(n1), .ZN(n133) );
  XNOR2_X1 U9 ( .A(n117), .B(n140), .ZN(result[22]) );
  INV_X1 U10 ( .A(n101), .ZN(n29) );
  AOI22_X1 U11 ( .A1(b[26]), .A2(a[26]), .B1(n7), .B2(n144), .ZN(n122) );
  AOI22_X1 U12 ( .A1(b[13]), .A2(a[13]), .B1(n21), .B2(n130), .ZN(n109) );
  OAI22_X1 U13 ( .A1(n11), .A2(n2), .B1(n150), .B2(n151), .ZN(cout) );
  INV_X1 U14 ( .A(n118), .ZN(n10) );
  INV_X1 U15 ( .A(n123), .ZN(n5) );
  AOI22_X1 U16 ( .A1(b[25]), .A2(a[25]), .B1(n8), .B2(n143), .ZN(n121) );
  INV_X1 U17 ( .A(n111), .ZN(n18) );
  INV_X1 U18 ( .A(n115), .ZN(n14) );
  INV_X1 U19 ( .A(n105), .ZN(n24) );
  AOI22_X1 U20 ( .A1(b[7]), .A2(a[7]), .B1(n27), .B2(n156), .ZN(n104) );
  INV_X1 U21 ( .A(n109), .ZN(n20) );
  INV_X1 U22 ( .A(n124), .ZN(n4) );
  AOI22_X1 U23 ( .A1(b[16]), .A2(a[16]), .B1(n18), .B2(n133), .ZN(n112) );
  AOI22_X1 U24 ( .A1(b[19]), .A2(a[19]), .B1(n15), .B2(n136), .ZN(n115) );
  INV_X1 U25 ( .A(n121), .ZN(n7) );
  AOI22_X1 U26 ( .A1(b[24]), .A2(a[24]), .B1(n9), .B2(n142), .ZN(n120) );
  AOI22_X1 U27 ( .A1(b[6]), .A2(a[6]), .B1(n28), .B2(n155), .ZN(n103) );
  AOI22_X1 U28 ( .A1(b[28]), .A2(a[28]), .B1(n5), .B2(n146), .ZN(n124) );
  AOI22_X1 U29 ( .A1(b[29]), .A2(a[29]), .B1(n4), .B2(n147), .ZN(n125) );
  AOI22_X1 U30 ( .A1(b[10]), .A2(a[10]), .B1(n24), .B2(n127), .ZN(n106) );
  AOI22_X1 U31 ( .A1(b[18]), .A2(a[18]), .B1(n16), .B2(n135), .ZN(n114) );
  AOI22_X1 U32 ( .A1(b[4]), .A2(a[4]), .B1(n30), .B2(n153), .ZN(n101) );
  AOI22_X1 U33 ( .A1(b[22]), .A2(a[22]), .B1(n12), .B2(n140), .ZN(n118) );
  AOI22_X1 U34 ( .A1(b[14]), .A2(a[14]), .B1(n20), .B2(n131), .ZN(n110) );
  INV_X1 U35 ( .A(n107), .ZN(n22) );
  AOI22_X1 U36 ( .A1(b[9]), .A2(a[9]), .B1(n25), .B2(n159), .ZN(n105) );
  AOI22_X1 U37 ( .A1(b[21]), .A2(a[21]), .B1(n13), .B2(n139), .ZN(n117) );
  AOI22_X1 U38 ( .A1(b[30]), .A2(a[30]), .B1(n3), .B2(n149), .ZN(n150) );
  AOI22_X1 U39 ( .A1(b[20]), .A2(a[20]), .B1(n14), .B2(n138), .ZN(n116) );
  INV_X1 U40 ( .A(n125), .ZN(n3) );
  AOI22_X1 U41 ( .A1(b[8]), .A2(a[8]), .B1(n26), .B2(n157), .ZN(n158) );
  INV_X1 U42 ( .A(n120), .ZN(n8) );
  INV_X1 U43 ( .A(n119), .ZN(n9) );
  INV_X1 U44 ( .A(n114), .ZN(n15) );
  INV_X1 U45 ( .A(n113), .ZN(n16) );
  INV_X1 U46 ( .A(n110), .ZN(n19) );
  INV_X1 U47 ( .A(n108), .ZN(n21) );
  INV_X1 U48 ( .A(n104), .ZN(n26) );
  INV_X1 U49 ( .A(n102), .ZN(n28) );
  INV_X1 U50 ( .A(n99), .ZN(n31) );
  AOI22_X1 U51 ( .A1(b[2]), .A2(a[2]), .B1(n32), .B2(n148), .ZN(n99) );
  AOI22_X1 U52 ( .A1(b[11]), .A2(a[11]), .B1(n23), .B2(n128), .ZN(n107) );
  AOI22_X1 U53 ( .A1(b[15]), .A2(a[15]), .B1(n19), .B2(n132), .ZN(n111) );
  AOI22_X1 U54 ( .A1(b[12]), .A2(a[12]), .B1(n22), .B2(n129), .ZN(n108) );
  AOI22_X1 U55 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(n152), .ZN(n100) );
  AOI22_X1 U56 ( .A1(b[5]), .A2(a[5]), .B1(n29), .B2(n154), .ZN(n102) );
  AOI22_X1 U57 ( .A1(b[23]), .A2(a[23]), .B1(n10), .B2(n141), .ZN(n119) );
  AOI22_X1 U58 ( .A1(b[17]), .A2(a[17]), .B1(n17), .B2(n134), .ZN(n113) );
  INV_X1 U59 ( .A(n122), .ZN(n6) );
  INV_X1 U60 ( .A(n117), .ZN(n12) );
  INV_X1 U61 ( .A(n116), .ZN(n13) );
  INV_X1 U62 ( .A(n112), .ZN(n17) );
  INV_X1 U63 ( .A(n106), .ZN(n23) );
  XNOR2_X1 U64 ( .A(n159), .B(n158), .ZN(result[9]) );
  INV_X1 U65 ( .A(n158), .ZN(n25) );
  INV_X1 U82 ( .A(n103), .ZN(n27) );
  AOI22_X1 U112 ( .A1(b[1]), .A2(a[1]), .B1(n96), .B2(n137), .ZN(n98) );
  AOI22_X1 U129 ( .A1(b[27]), .A2(a[27]), .B1(n6), .B2(n145), .ZN(n123) );
endmodule


module carryLookAheadAdder_20 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n12), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n13), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n14), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n15), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n16), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n17), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  AOI22_X1 U1 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  INV_X1 U2 ( .A(a[31]), .ZN(n1) );
  OAI22_X1 U3 ( .A1(n11), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U4 ( .A(b[31]), .ZN(n11) );
  INV_X1 U5 ( .A(n103), .ZN(n25) );
  INV_X1 U6 ( .A(n99), .ZN(n29) );
  INV_X1 U7 ( .A(n96), .ZN(n32) );
  AOI22_X1 U8 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  AOI22_X1 U9 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  INV_X1 U10 ( .A(n107), .ZN(n20) );
  AOI22_X1 U11 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  INV_X1 U12 ( .A(n98), .ZN(n30) );
  INV_X1 U13 ( .A(n118), .ZN(n8) );
  INV_X1 U14 ( .A(n117), .ZN(n9) );
  XNOR2_X1 U15 ( .A(n124), .B(n148), .ZN(result[30]) );
  AOI22_X1 U16 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  INV_X1 U17 ( .A(n104), .ZN(n23) );
  AOI22_X1 U18 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  INV_X1 U19 ( .A(n100), .ZN(n28) );
  INV_X1 U20 ( .A(n120), .ZN(n6) );
  INV_X1 U21 ( .A(n116), .ZN(n10) );
  AOI22_X1 U22 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  INV_X1 U23 ( .A(n106), .ZN(n21) );
  AOI22_X1 U24 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  INV_X1 U25 ( .A(n101), .ZN(n27) );
  INV_X1 U26 ( .A(n97), .ZN(n31) );
  AOI22_X1 U27 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  AOI22_X1 U28 ( .A1(b[18]), .A2(a[18]), .B1(n15), .B2(n134), .ZN(n113) );
  AOI22_X1 U29 ( .A1(b[17]), .A2(a[17]), .B1(n16), .B2(n133), .ZN(n112) );
  AOI22_X1 U30 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  AOI22_X1 U31 ( .A1(b[21]), .A2(a[21]), .B1(n12), .B2(n138), .ZN(n116) );
  AOI22_X1 U32 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  INV_X1 U33 ( .A(n124), .ZN(n2) );
  INV_X1 U34 ( .A(n122), .ZN(n4) );
  INV_X1 U35 ( .A(n114), .ZN(n13) );
  INV_X1 U36 ( .A(n112), .ZN(n15) );
  AOI22_X1 U37 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
  AOI22_X1 U38 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  AOI22_X1 U39 ( .A1(b[20]), .A2(a[20]), .B1(n13), .B2(n137), .ZN(n115) );
  AOI22_X1 U40 ( .A1(b[19]), .A2(a[19]), .B1(n14), .B2(n135), .ZN(n114) );
  AOI22_X1 U41 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U42 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  INV_X1 U43 ( .A(n108), .ZN(n19) );
  INV_X1 U44 ( .A(n110), .ZN(n17) );
  AOI22_X1 U45 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  AOI22_X1 U46 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  INV_X1 U47 ( .A(n123), .ZN(n3) );
  AOI22_X1 U48 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U49 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U50 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U51 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U52 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  AOI22_X1 U53 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  INV_X1 U54 ( .A(n121), .ZN(n5) );
  INV_X1 U55 ( .A(n119), .ZN(n7) );
  INV_X1 U56 ( .A(n115), .ZN(n12) );
  INV_X1 U57 ( .A(n113), .ZN(n14) );
  INV_X1 U58 ( .A(n111), .ZN(n16) );
  INV_X1 U59 ( .A(n109), .ZN(n18) );
  INV_X1 U60 ( .A(n105), .ZN(n22) );
  XNOR2_X1 U61 ( .A(n158), .B(n157), .ZN(result[9]) );
  INV_X1 U62 ( .A(n157), .ZN(n24) );
  AOI22_X1 U63 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  INV_X1 U64 ( .A(n102), .ZN(n26) );
  AOI22_X1 U65 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U73 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
endmodule


module carryLookAheadAdder_19 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n13), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n14), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n15), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n16), .Z(result[17]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  OAI22_X1 U1 ( .A1(n12), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U2 ( .A(b[31]), .ZN(n12) );
  INV_X1 U3 ( .A(a[31]), .ZN(n1) );
  INV_X1 U4 ( .A(n124), .ZN(n2) );
  INV_X1 U5 ( .A(n116), .ZN(n10) );
  INV_X1 U6 ( .A(n101), .ZN(n27) );
  INV_X1 U7 ( .A(n99), .ZN(n29) );
  INV_X1 U8 ( .A(n97), .ZN(n31) );
  INV_X1 U9 ( .A(n96), .ZN(n32) );
  AOI22_X1 U10 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  AOI22_X1 U11 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  INV_X1 U12 ( .A(n98), .ZN(n30) );
  INV_X1 U13 ( .A(n121), .ZN(n5) );
  INV_X1 U14 ( .A(n114), .ZN(n13) );
  XNOR2_X1 U15 ( .A(n110), .B(n132), .ZN(result[16]) );
  AOI22_X1 U16 ( .A1(b[20]), .A2(a[20]), .B1(n13), .B2(n137), .ZN(n115) );
  INV_X1 U17 ( .A(n103), .ZN(n25) );
  INV_X1 U18 ( .A(n105), .ZN(n22) );
  INV_X1 U19 ( .A(n110), .ZN(n17) );
  INV_X1 U20 ( .A(n120), .ZN(n6) );
  INV_X1 U21 ( .A(n108), .ZN(n19) );
  AOI22_X1 U22 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  INV_X1 U23 ( .A(n113), .ZN(n14) );
  INV_X1 U24 ( .A(n117), .ZN(n9) );
  AOI22_X1 U25 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  AOI22_X1 U26 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  AOI22_X1 U27 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  INV_X1 U28 ( .A(n102), .ZN(n26) );
  AOI22_X1 U29 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U30 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U31 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U32 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
  INV_X1 U33 ( .A(n107), .ZN(n20) );
  AOI22_X1 U34 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  AOI22_X1 U35 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  AOI22_X1 U36 ( .A1(b[19]), .A2(a[19]), .B1(n14), .B2(n135), .ZN(n114) );
  AOI22_X1 U37 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U38 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  AOI22_X1 U39 ( .A1(b[18]), .A2(a[18]), .B1(n15), .B2(n134), .ZN(n113) );
  AOI22_X1 U40 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U41 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  INV_X1 U42 ( .A(n123), .ZN(n3) );
  INV_X1 U43 ( .A(n122), .ZN(n4) );
  INV_X1 U44 ( .A(n119), .ZN(n7) );
  INV_X1 U45 ( .A(n118), .ZN(n8) );
  INV_X1 U46 ( .A(n115), .ZN(n11) );
  INV_X1 U47 ( .A(n112), .ZN(n15) );
  INV_X1 U48 ( .A(n111), .ZN(n16) );
  AOI22_X1 U49 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  AOI22_X1 U50 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  AOI22_X1 U51 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U52 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U53 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  AOI22_X1 U54 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U55 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  INV_X1 U56 ( .A(n109), .ZN(n18) );
  INV_X1 U57 ( .A(n106), .ZN(n21) );
  INV_X1 U58 ( .A(n104), .ZN(n23) );
  XNOR2_X1 U59 ( .A(n158), .B(n157), .ZN(result[9]) );
  INV_X1 U60 ( .A(n157), .ZN(n24) );
  INV_X1 U61 ( .A(n100), .ZN(n28) );
  AOI22_X1 U62 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U63 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  AOI22_X1 U64 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  AOI22_X1 U65 ( .A1(b[17]), .A2(a[17]), .B1(n16), .B2(n133), .ZN(n112) );
  AOI22_X1 U89 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
endmodule


module carryLookAheadAdder_18 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n14), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n15), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n16), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n17), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  INV_X1 U1 ( .A(a[31]), .ZN(n1) );
  OAI22_X1 U2 ( .A1(n13), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U3 ( .A(b[31]), .ZN(n13) );
  INV_X1 U4 ( .A(n115), .ZN(n11) );
  INV_X1 U5 ( .A(n99), .ZN(n29) );
  INV_X1 U6 ( .A(n97), .ZN(n31) );
  INV_X1 U7 ( .A(n96), .ZN(n32) );
  AOI22_X1 U8 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U9 ( .A(n98), .ZN(n30) );
  INV_X1 U10 ( .A(n103), .ZN(n25) );
  INV_X1 U11 ( .A(n100), .ZN(n28) );
  AOI22_X1 U12 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  INV_X1 U13 ( .A(n122), .ZN(n4) );
  INV_X1 U14 ( .A(n109), .ZN(n18) );
  AOI22_X1 U15 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  INV_X1 U16 ( .A(n106), .ZN(n21) );
  INV_X1 U17 ( .A(n120), .ZN(n6) );
  AOI22_X1 U18 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  AOI22_X1 U19 ( .A1(b[18]), .A2(a[18]), .B1(n15), .B2(n134), .ZN(n113) );
  INV_X1 U20 ( .A(n101), .ZN(n27) );
  INV_X1 U21 ( .A(n114), .ZN(n12) );
  INV_X1 U22 ( .A(n112), .ZN(n15) );
  INV_X1 U23 ( .A(n108), .ZN(n19) );
  INV_X1 U24 ( .A(n107), .ZN(n20) );
  AOI22_X1 U25 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U26 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U27 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U28 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  AOI22_X1 U29 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U30 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  AOI22_X1 U31 ( .A1(b[19]), .A2(a[19]), .B1(n14), .B2(n135), .ZN(n114) );
  INV_X1 U32 ( .A(n118), .ZN(n8) );
  INV_X1 U33 ( .A(n117), .ZN(n9) );
  INV_X1 U34 ( .A(n116), .ZN(n10) );
  INV_X1 U35 ( .A(n111), .ZN(n16) );
  AOI22_X1 U36 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  AOI22_X1 U37 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  AOI22_X1 U38 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  AOI22_X1 U39 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  INV_X1 U40 ( .A(n123), .ZN(n3) );
  INV_X1 U41 ( .A(n124), .ZN(n2) );
  AOI22_X1 U42 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U43 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  AOI22_X1 U44 ( .A1(b[17]), .A2(a[17]), .B1(n16), .B2(n133), .ZN(n112) );
  AOI22_X1 U45 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U46 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  AOI22_X1 U47 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  AOI22_X1 U48 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  AOI22_X1 U49 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U50 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  AOI22_X1 U51 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  INV_X1 U52 ( .A(n110), .ZN(n17) );
  INV_X1 U53 ( .A(n105), .ZN(n22) );
  INV_X1 U54 ( .A(n104), .ZN(n23) );
  XNOR2_X1 U55 ( .A(n158), .B(n157), .ZN(result[9]) );
  INV_X1 U56 ( .A(n157), .ZN(n24) );
  INV_X1 U57 ( .A(n102), .ZN(n26) );
  AOI22_X1 U58 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  INV_X1 U59 ( .A(n121), .ZN(n5) );
  INV_X1 U60 ( .A(n119), .ZN(n7) );
  INV_X1 U61 ( .A(n113), .ZN(n14) );
  AOI22_X1 U62 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
  AOI22_X1 U63 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U64 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  AOI22_X1 U65 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
endmodule


module carryLookAheadAdder_17 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n15), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n16), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n17), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  XOR2_X1 U1 ( .A(a[16]), .B(b[16]), .Z(n132) );
  AOI22_X1 U2 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  INV_X1 U3 ( .A(n124), .ZN(n2) );
  OAI22_X1 U4 ( .A1(n14), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U5 ( .A(b[31]), .ZN(n14) );
  INV_X1 U6 ( .A(a[31]), .ZN(n1) );
  INV_X1 U7 ( .A(n120), .ZN(n6) );
  INV_X1 U8 ( .A(n97), .ZN(n31) );
  INV_X1 U9 ( .A(n96), .ZN(n32) );
  AOI22_X1 U10 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U11 ( .A(n99), .ZN(n29) );
  INV_X1 U12 ( .A(n102), .ZN(n26) );
  INV_X1 U13 ( .A(n103), .ZN(n25) );
  INV_X1 U14 ( .A(n114), .ZN(n12) );
  INV_X1 U15 ( .A(n107), .ZN(n20) );
  AOI22_X1 U16 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  INV_X1 U17 ( .A(n109), .ZN(n18) );
  INV_X1 U18 ( .A(n113), .ZN(n13) );
  INV_X1 U19 ( .A(n118), .ZN(n8) );
  INV_X1 U20 ( .A(n101), .ZN(n27) );
  INV_X1 U21 ( .A(n121), .ZN(n5) );
  INV_X1 U22 ( .A(n116), .ZN(n10) );
  INV_X1 U23 ( .A(n115), .ZN(n11) );
  INV_X1 U24 ( .A(n111), .ZN(n16) );
  INV_X1 U25 ( .A(n110), .ZN(n17) );
  INV_X1 U26 ( .A(n106), .ZN(n21) );
  INV_X1 U27 ( .A(n104), .ZN(n23) );
  INV_X1 U28 ( .A(n100), .ZN(n28) );
  AOI22_X1 U29 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  INV_X1 U30 ( .A(n105), .ZN(n22) );
  AOI22_X1 U31 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U32 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  AOI22_X1 U33 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  AOI22_X1 U34 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  AOI22_X1 U35 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  INV_X1 U36 ( .A(n123), .ZN(n3) );
  AOI22_X1 U37 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  AOI22_X1 U38 ( .A1(b[18]), .A2(a[18]), .B1(n15), .B2(n134), .ZN(n113) );
  AOI22_X1 U39 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U40 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U41 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U42 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  AOI22_X1 U43 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  AOI22_X1 U44 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U45 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U46 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U47 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U48 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U49 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  INV_X1 U50 ( .A(n122), .ZN(n4) );
  INV_X1 U51 ( .A(n119), .ZN(n7) );
  INV_X1 U52 ( .A(n117), .ZN(n9) );
  INV_X1 U53 ( .A(n112), .ZN(n15) );
  AOI22_X1 U54 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
  AOI22_X1 U55 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  INV_X1 U56 ( .A(n108), .ZN(n19) );
  XNOR2_X1 U57 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U58 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  INV_X1 U59 ( .A(n157), .ZN(n24) );
  INV_X1 U60 ( .A(n98), .ZN(n30) );
  AOI22_X1 U61 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U62 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U63 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  AOI22_X1 U64 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  AOI22_X1 U65 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  AOI22_X1 U112 ( .A1(b[17]), .A2(a[17]), .B1(n16), .B2(n133), .ZN(n112) );
endmodule


module carryLookAheadAdder_16 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n16), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n17), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  INV_X1 U1 ( .A(a[31]), .ZN(n1) );
  INV_X1 U2 ( .A(n123), .ZN(n3) );
  INV_X1 U3 ( .A(n117), .ZN(n9) );
  INV_X1 U4 ( .A(n122), .ZN(n4) );
  OAI22_X1 U5 ( .A1(n15), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U6 ( .A(b[31]), .ZN(n15) );
  INV_X1 U7 ( .A(n96), .ZN(n32) );
  AOI22_X1 U8 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U9 ( .A(n100), .ZN(n28) );
  INV_X1 U10 ( .A(n99), .ZN(n29) );
  AOI22_X1 U11 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  AOI22_X1 U12 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  INV_X1 U13 ( .A(n121), .ZN(n5) );
  XNOR2_X1 U14 ( .A(n106), .B(n128), .ZN(result[12]) );
  INV_X1 U15 ( .A(n111), .ZN(n16) );
  INV_X1 U16 ( .A(n157), .ZN(n24) );
  INV_X1 U17 ( .A(n98), .ZN(n30) );
  INV_X1 U18 ( .A(n97), .ZN(n31) );
  XNOR2_X1 U19 ( .A(n108), .B(n130), .ZN(result[14]) );
  INV_X1 U20 ( .A(n116), .ZN(n10) );
  INV_X1 U21 ( .A(n104), .ZN(n23) );
  INV_X1 U22 ( .A(n105), .ZN(n22) );
  INV_X1 U23 ( .A(n113), .ZN(n13) );
  INV_X1 U24 ( .A(n110), .ZN(n17) );
  INV_X1 U25 ( .A(n108), .ZN(n19) );
  INV_X1 U26 ( .A(n120), .ZN(n6) );
  INV_X1 U27 ( .A(n124), .ZN(n2) );
  AOI22_X1 U28 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  AOI22_X1 U29 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  INV_X1 U30 ( .A(n101), .ZN(n27) );
  AOI22_X1 U31 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U32 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  AOI22_X1 U33 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  AOI22_X1 U34 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
  AOI22_X1 U35 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  AOI22_X1 U36 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U37 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U38 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  AOI22_X1 U39 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  INV_X1 U40 ( .A(n114), .ZN(n12) );
  INV_X1 U41 ( .A(n112), .ZN(n14) );
  INV_X1 U42 ( .A(n107), .ZN(n20) );
  INV_X1 U43 ( .A(n106), .ZN(n21) );
  INV_X1 U44 ( .A(n103), .ZN(n25) );
  INV_X1 U45 ( .A(n102), .ZN(n26) );
  AOI22_X1 U46 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U47 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  AOI22_X1 U48 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U49 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U50 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U51 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U52 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U53 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U54 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U55 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  AOI22_X1 U56 ( .A1(b[17]), .A2(a[17]), .B1(n16), .B2(n133), .ZN(n112) );
  INV_X1 U57 ( .A(n119), .ZN(n7) );
  INV_X1 U58 ( .A(n118), .ZN(n8) );
  AOI22_X1 U59 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  INV_X1 U60 ( .A(n115), .ZN(n11) );
  INV_X1 U61 ( .A(n109), .ZN(n18) );
  AOI22_X1 U62 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  AOI22_X1 U63 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  AOI22_X1 U64 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  XNOR2_X1 U65 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U91 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  AOI22_X1 U93 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
endmodule


module carryLookAheadAdder_15 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  XOR2_X1 U1 ( .A(a[11]), .B(b[11]), .Z(n127) );
  INV_X1 U2 ( .A(b[31]), .ZN(n16) );
  INV_X1 U3 ( .A(n122), .ZN(n4) );
  INV_X1 U4 ( .A(n120), .ZN(n6) );
  INV_X1 U5 ( .A(n124), .ZN(n2) );
  AOI22_X1 U6 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  INV_X1 U7 ( .A(a[31]), .ZN(n1) );
  INV_X1 U8 ( .A(n97), .ZN(n31) );
  INV_X1 U9 ( .A(n96), .ZN(n32) );
  AOI22_X1 U10 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U11 ( .A(n101), .ZN(n27) );
  INV_X1 U12 ( .A(n99), .ZN(n29) );
  INV_X1 U13 ( .A(n103), .ZN(n25) );
  XNOR2_X1 U14 ( .A(n110), .B(n132), .ZN(result[16]) );
  INV_X1 U15 ( .A(n107), .ZN(n20) );
  INV_X1 U16 ( .A(n117), .ZN(n9) );
  INV_X1 U17 ( .A(n116), .ZN(n10) );
  INV_X1 U18 ( .A(n113), .ZN(n13) );
  INV_X1 U19 ( .A(n114), .ZN(n12) );
  AOI22_X1 U20 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  OAI22_X1 U21 ( .A1(n16), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U22 ( .A(n123), .ZN(n3) );
  AOI22_X1 U23 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  INV_X1 U24 ( .A(n108), .ZN(n19) );
  INV_X1 U25 ( .A(n106), .ZN(n21) );
  AOI22_X1 U26 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  AOI22_X1 U27 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  INV_X1 U28 ( .A(n105), .ZN(n22) );
  AOI22_X1 U29 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  AOI22_X1 U30 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U31 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  AOI22_X1 U32 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  INV_X1 U33 ( .A(n102), .ZN(n26) );
  AOI22_X1 U34 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U35 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  INV_X1 U36 ( .A(n115), .ZN(n11) );
  AOI22_X1 U37 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U38 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  AOI22_X1 U39 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  AOI22_X1 U40 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U41 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  AOI22_X1 U42 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U43 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  AOI22_X1 U44 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U45 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U46 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U47 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U48 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U49 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  INV_X1 U50 ( .A(n121), .ZN(n5) );
  INV_X1 U51 ( .A(n119), .ZN(n7) );
  INV_X1 U52 ( .A(n118), .ZN(n8) );
  INV_X1 U53 ( .A(n112), .ZN(n14) );
  INV_X1 U54 ( .A(n111), .ZN(n15) );
  INV_X1 U55 ( .A(n110), .ZN(n17) );
  INV_X1 U56 ( .A(n109), .ZN(n18) );
  INV_X1 U57 ( .A(n104), .ZN(n23) );
  INV_X1 U58 ( .A(n157), .ZN(n24) );
  INV_X1 U59 ( .A(n100), .ZN(n28) );
  INV_X1 U60 ( .A(n98), .ZN(n30) );
  AOI22_X1 U61 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U62 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
  AOI22_X1 U63 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  AOI22_X1 U64 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  XNOR2_X1 U65 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U89 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  AOI22_X1 U117 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
endmodule


module carryLookAheadAdder_14 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  XOR2_X1 U1 ( .A(a[11]), .B(b[11]), .Z(n127) );
  AOI22_X1 U2 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  INV_X1 U3 ( .A(a[31]), .ZN(n1) );
  INV_X1 U4 ( .A(n124), .ZN(n2) );
  OAI22_X1 U5 ( .A1(n17), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U6 ( .A(b[31]), .ZN(n17) );
  INV_X1 U7 ( .A(n120), .ZN(n6) );
  INV_X1 U8 ( .A(n122), .ZN(n4) );
  INV_X1 U9 ( .A(n96), .ZN(n32) );
  AOI22_X1 U10 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U11 ( .A(n99), .ZN(n29) );
  INV_X1 U12 ( .A(n97), .ZN(n31) );
  INV_X1 U13 ( .A(n110), .ZN(n16) );
  INV_X1 U14 ( .A(n101), .ZN(n27) );
  INV_X1 U15 ( .A(n102), .ZN(n26) );
  INV_X1 U16 ( .A(n118), .ZN(n8) );
  INV_X1 U17 ( .A(n112), .ZN(n14) );
  XNOR2_X1 U18 ( .A(n127), .B(n105), .ZN(result[11]) );
  INV_X1 U19 ( .A(n106), .ZN(n21) );
  INV_X1 U20 ( .A(n103), .ZN(n25) );
  INV_X1 U21 ( .A(n98), .ZN(n30) );
  INV_X1 U22 ( .A(n111), .ZN(n15) );
  INV_X1 U23 ( .A(n114), .ZN(n12) );
  INV_X1 U24 ( .A(n117), .ZN(n9) );
  INV_X1 U25 ( .A(n108), .ZN(n19) );
  AOI22_X1 U26 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  AOI22_X1 U27 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  INV_X1 U28 ( .A(n123), .ZN(n3) );
  AOI22_X1 U29 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  AOI22_X1 U30 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n132), .ZN(n111) );
  INV_X1 U31 ( .A(n104), .ZN(n23) );
  AOI22_X1 U32 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  AOI22_X1 U33 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U34 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  AOI22_X1 U35 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  AOI22_X1 U36 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U37 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  AOI22_X1 U38 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  AOI22_X1 U39 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  AOI22_X1 U40 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  AOI22_X1 U41 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  AOI22_X1 U42 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U43 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U44 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  AOI22_X1 U45 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U46 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U47 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U48 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U49 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U50 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U51 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U52 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  AOI22_X1 U53 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  INV_X1 U54 ( .A(n121), .ZN(n5) );
  INV_X1 U55 ( .A(n119), .ZN(n7) );
  INV_X1 U56 ( .A(n116), .ZN(n10) );
  INV_X1 U57 ( .A(n115), .ZN(n11) );
  INV_X1 U58 ( .A(n113), .ZN(n13) );
  INV_X1 U59 ( .A(n109), .ZN(n18) );
  INV_X1 U60 ( .A(n107), .ZN(n20) );
  INV_X1 U61 ( .A(n105), .ZN(n22) );
  XNOR2_X1 U62 ( .A(n158), .B(n157), .ZN(result[9]) );
  INV_X1 U63 ( .A(n157), .ZN(n24) );
  INV_X1 U64 ( .A(n100), .ZN(n28) );
  AOI22_X1 U65 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U94 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  AOI22_X1 U117 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
endmodule


module carryLookAheadAdder_13 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n17), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n20), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  XOR2_X1 U1 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U2 ( .A(a[9]), .B(b[9]), .Z(n158) );
  AOI22_X1 U3 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  INV_X1 U4 ( .A(n124), .ZN(n2) );
  INV_X1 U5 ( .A(a[31]), .ZN(n1) );
  INV_X1 U6 ( .A(n123), .ZN(n3) );
  INV_X1 U7 ( .A(n118), .ZN(n8) );
  INV_X1 U8 ( .A(n122), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n18), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U10 ( .A(b[31]), .ZN(n18) );
  INV_X1 U11 ( .A(n96), .ZN(n32) );
  AOI22_X1 U12 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  AOI22_X1 U13 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  INV_X1 U14 ( .A(n97), .ZN(n31) );
  INV_X1 U15 ( .A(n98), .ZN(n30) );
  INV_X1 U16 ( .A(n99), .ZN(n29) );
  AOI22_X1 U17 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  INV_X1 U18 ( .A(n108), .ZN(n19) );
  INV_X1 U19 ( .A(n109), .ZN(n17) );
  INV_X1 U20 ( .A(n103), .ZN(n25) );
  INV_X1 U21 ( .A(n102), .ZN(n26) );
  INV_X1 U22 ( .A(n113), .ZN(n13) );
  INV_X1 U23 ( .A(n107), .ZN(n20) );
  INV_X1 U24 ( .A(n115), .ZN(n11) );
  INV_X1 U25 ( .A(n117), .ZN(n9) );
  INV_X1 U26 ( .A(n101), .ZN(n27) );
  INV_X1 U27 ( .A(n112), .ZN(n14) );
  INV_X1 U28 ( .A(n110), .ZN(n16) );
  AOI22_X1 U29 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  AOI22_X1 U30 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  INV_X1 U31 ( .A(n111), .ZN(n15) );
  AOI22_X1 U32 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U33 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U34 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  AOI22_X1 U35 ( .A1(b[15]), .A2(a[15]), .B1(n17), .B2(n131), .ZN(n110) );
  AOI22_X1 U36 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  AOI22_X1 U37 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  AOI22_X1 U38 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  AOI22_X1 U39 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U40 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  AOI22_X1 U41 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U42 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  AOI22_X1 U43 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  INV_X1 U44 ( .A(n121), .ZN(n5) );
  INV_X1 U45 ( .A(n120), .ZN(n6) );
  AOI22_X1 U46 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U47 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  AOI22_X1 U48 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n132), .ZN(n111) );
  INV_X1 U49 ( .A(n119), .ZN(n7) );
  INV_X1 U50 ( .A(n116), .ZN(n10) );
  INV_X1 U51 ( .A(n114), .ZN(n12) );
  INV_X1 U52 ( .A(n106), .ZN(n21) );
  INV_X1 U53 ( .A(n105), .ZN(n22) );
  INV_X1 U54 ( .A(n104), .ZN(n23) );
  XNOR2_X1 U55 ( .A(n158), .B(n157), .ZN(result[9]) );
  INV_X1 U56 ( .A(n157), .ZN(n24) );
  INV_X1 U57 ( .A(n100), .ZN(n28) );
  AOI22_X1 U58 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U59 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U60 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  AOI22_X1 U61 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  AOI22_X1 U62 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  AOI22_X1 U63 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U64 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  AOI22_X1 U65 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  AOI22_X1 U117 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U119 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
endmodule


module carryLookAheadAdder_12 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n26), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n27), .Z(result[7]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n3), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n4), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n5), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n6), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n7), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n8), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n9), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n10), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n11), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n12), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n13), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n14), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n15), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n16), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n17), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n18), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n19), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n21), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n22), .B(n128), .Z(result[12]) );
  XOR2_X1 U95 ( .A(n24), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n2), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  XNOR2_X1 U1 ( .A(n101), .B(n154), .ZN(result[6]) );
  XOR2_X1 U2 ( .A(a[5]), .B(b[5]), .Z(n153) );
  AOI22_X1 U3 ( .A1(b[30]), .A2(a[30]), .B1(n3), .B2(n148), .ZN(n149) );
  INV_X1 U4 ( .A(b[31]), .ZN(n20) );
  INV_X1 U5 ( .A(n118), .ZN(n9) );
  INV_X1 U6 ( .A(n120), .ZN(n7) );
  INV_X1 U7 ( .A(n122), .ZN(n5) );
  INV_X1 U8 ( .A(n106), .ZN(n22) );
  INV_X1 U9 ( .A(a[31]), .ZN(n2) );
  INV_X1 U10 ( .A(n96), .ZN(n32) );
  AOI22_X1 U11 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U12 ( .A(n97), .ZN(n31) );
  INV_X1 U13 ( .A(n101), .ZN(n1) );
  INV_X1 U14 ( .A(n114), .ZN(n13) );
  XNOR2_X1 U15 ( .A(n127), .B(n105), .ZN(result[11]) );
  INV_X1 U16 ( .A(n105), .ZN(n23) );
  INV_X1 U17 ( .A(n100), .ZN(n28) );
  INV_X1 U18 ( .A(n115), .ZN(n12) );
  INV_X1 U19 ( .A(n102), .ZN(n27) );
  INV_X1 U20 ( .A(n104), .ZN(n24) );
  AOI22_X1 U21 ( .A1(b[11]), .A2(a[11]), .B1(n23), .B2(n127), .ZN(n106) );
  INV_X1 U22 ( .A(n112), .ZN(n15) );
  INV_X1 U23 ( .A(n110), .ZN(n17) );
  INV_X1 U24 ( .A(n108), .ZN(n19) );
  INV_X1 U25 ( .A(n103), .ZN(n26) );
  INV_X1 U26 ( .A(n99), .ZN(n29) );
  INV_X1 U27 ( .A(n98), .ZN(n30) );
  AOI22_X1 U28 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U29 ( .A1(b[29]), .A2(a[29]), .B1(n4), .B2(n146), .ZN(n124) );
  AOI22_X1 U30 ( .A1(b[14]), .A2(a[14]), .B1(n19), .B2(n130), .ZN(n109) );
  AOI22_X1 U31 ( .A1(b[20]), .A2(a[20]), .B1(n13), .B2(n137), .ZN(n115) );
  AOI22_X1 U32 ( .A1(b[9]), .A2(a[9]), .B1(n25), .B2(n158), .ZN(n104) );
  INV_X1 U33 ( .A(n124), .ZN(n3) );
  INV_X1 U34 ( .A(n123), .ZN(n4) );
  AOI22_X1 U35 ( .A1(b[24]), .A2(a[24]), .B1(n9), .B2(n141), .ZN(n119) );
  AOI22_X1 U36 ( .A1(b[22]), .A2(a[22]), .B1(n11), .B2(n139), .ZN(n117) );
  AOI22_X1 U37 ( .A1(b[6]), .A2(a[6]), .B1(n1), .B2(n154), .ZN(n102) );
  AOI22_X1 U38 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U39 ( .A1(b[13]), .A2(a[13]), .B1(n21), .B2(n129), .ZN(n108) );
  AOI22_X1 U40 ( .A1(b[25]), .A2(a[25]), .B1(n8), .B2(n142), .ZN(n120) );
  AOI22_X1 U41 ( .A1(b[18]), .A2(a[18]), .B1(n15), .B2(n134), .ZN(n113) );
  AOI22_X1 U42 ( .A1(b[27]), .A2(a[27]), .B1(n6), .B2(n144), .ZN(n122) );
  AOI22_X1 U43 ( .A1(b[23]), .A2(a[23]), .B1(n10), .B2(n140), .ZN(n118) );
  AOI22_X1 U44 ( .A1(b[12]), .A2(a[12]), .B1(n22), .B2(n128), .ZN(n107) );
  AOI22_X1 U45 ( .A1(b[17]), .A2(a[17]), .B1(n16), .B2(n133), .ZN(n112) );
  AOI22_X1 U46 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U47 ( .A1(b[19]), .A2(a[19]), .B1(n14), .B2(n135), .ZN(n114) );
  INV_X1 U48 ( .A(n116), .ZN(n11) );
  AOI22_X1 U49 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U50 ( .A1(b[8]), .A2(a[8]), .B1(n26), .B2(n156), .ZN(n157) );
  AOI22_X1 U51 ( .A1(b[21]), .A2(a[21]), .B1(n12), .B2(n138), .ZN(n116) );
  AOI22_X1 U52 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U53 ( .A1(b[15]), .A2(a[15]), .B1(n18), .B2(n131), .ZN(n110) );
  AOI22_X1 U54 ( .A1(b[28]), .A2(a[28]), .B1(n5), .B2(n145), .ZN(n123) );
  AOI22_X1 U55 ( .A1(b[16]), .A2(a[16]), .B1(n17), .B2(n132), .ZN(n111) );
  AOI22_X1 U56 ( .A1(b[26]), .A2(a[26]), .B1(n7), .B2(n143), .ZN(n121) );
  OAI22_X1 U57 ( .A1(n20), .A2(n2), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U58 ( .A(n121), .ZN(n6) );
  INV_X1 U59 ( .A(n119), .ZN(n8) );
  INV_X1 U60 ( .A(n117), .ZN(n10) );
  INV_X1 U61 ( .A(n113), .ZN(n14) );
  INV_X1 U62 ( .A(n111), .ZN(n16) );
  INV_X1 U63 ( .A(n109), .ZN(n18) );
  INV_X1 U64 ( .A(n107), .ZN(n21) );
  XNOR2_X1 U65 ( .A(n158), .B(n157), .ZN(result[9]) );
  INV_X1 U68 ( .A(n157), .ZN(n25) );
  AOI22_X1 U94 ( .A1(b[7]), .A2(a[7]), .B1(n27), .B2(n155), .ZN(n103) );
  AOI22_X1 U123 ( .A1(b[10]), .A2(a[10]), .B1(n24), .B2(n126), .ZN(n105) );
endmodule


module carryLookAheadAdder_11 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n26), .B(n155), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n28), .B(n153), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n17), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n18), .B(n130), .Z(result[14]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  XOR2_X1 U1 ( .A(a[9]), .B(b[9]), .Z(n158) );
  INV_X1 U2 ( .A(b[31]), .ZN(n19) );
  INV_X1 U3 ( .A(a[31]), .ZN(n1) );
  INV_X1 U4 ( .A(n116), .ZN(n10) );
  INV_X1 U5 ( .A(n124), .ZN(n2) );
  AOI22_X1 U6 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U7 ( .A(n96), .ZN(n32) );
  AOI22_X1 U8 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  INV_X1 U9 ( .A(n99), .ZN(n29) );
  INV_X1 U10 ( .A(n98), .ZN(n30) );
  INV_X1 U11 ( .A(n115), .ZN(n11) );
  INV_X1 U12 ( .A(n97), .ZN(n31) );
  XNOR2_X1 U13 ( .A(n104), .B(n126), .ZN(result[10]) );
  XNOR2_X1 U14 ( .A(n129), .B(n107), .ZN(result[13]) );
  XNOR2_X1 U15 ( .A(n127), .B(n105), .ZN(result[11]) );
  INV_X1 U16 ( .A(n101), .ZN(n27) );
  INV_X1 U17 ( .A(n108), .ZN(n18) );
  INV_X1 U18 ( .A(n110), .ZN(n16) );
  INV_X1 U19 ( .A(n103), .ZN(n25) );
  INV_X1 U20 ( .A(n104), .ZN(n23) );
  AOI22_X1 U21 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  INV_X1 U22 ( .A(n106), .ZN(n21) );
  INV_X1 U23 ( .A(n100), .ZN(n28) );
  INV_X1 U24 ( .A(n120), .ZN(n6) );
  INV_X1 U25 ( .A(n118), .ZN(n8) );
  AOI22_X1 U26 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U27 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  AOI22_X1 U28 ( .A1(b[15]), .A2(a[15]), .B1(n17), .B2(n131), .ZN(n110) );
  AOI22_X1 U29 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  INV_X1 U30 ( .A(n122), .ZN(n4) );
  INV_X1 U31 ( .A(n121), .ZN(n5) );
  INV_X1 U32 ( .A(n114), .ZN(n12) );
  INV_X1 U33 ( .A(n111), .ZN(n15) );
  INV_X1 U34 ( .A(n105), .ZN(n22) );
  INV_X1 U35 ( .A(n102), .ZN(n26) );
  AOI22_X1 U36 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U37 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  AOI22_X1 U38 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U39 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  AOI22_X1 U40 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U41 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U42 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  AOI22_X1 U43 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U44 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U45 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U46 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  AOI22_X1 U47 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U48 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n132), .ZN(n111) );
  AOI22_X1 U49 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U50 ( .A1(b[14]), .A2(a[14]), .B1(n18), .B2(n130), .ZN(n109) );
  INV_X1 U51 ( .A(n123), .ZN(n3) );
  AOI22_X1 U52 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  AOI22_X1 U53 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  AOI22_X1 U54 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  AOI22_X1 U55 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U56 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  AOI22_X1 U57 ( .A1(b[13]), .A2(a[13]), .B1(n20), .B2(n129), .ZN(n108) );
  OAI22_X1 U58 ( .A1(n19), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U59 ( .A(n119), .ZN(n7) );
  INV_X1 U60 ( .A(n117), .ZN(n9) );
  INV_X1 U61 ( .A(n113), .ZN(n13) );
  INV_X1 U62 ( .A(n112), .ZN(n14) );
  INV_X1 U63 ( .A(n109), .ZN(n17) );
  INV_X1 U64 ( .A(n107), .ZN(n20) );
  XNOR2_X1 U65 ( .A(n158), .B(n157), .ZN(result[9]) );
  INV_X1 U92 ( .A(n157), .ZN(n24) );
  AOI22_X1 U94 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  AOI22_X1 U95 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  AOI22_X1 U119 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
endmodule


module carryLookAheadAdder_10 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n26), .B(n155), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n17), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n18), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n19), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n21), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  INV_X1 U1 ( .A(a[31]), .ZN(n1) );
  OAI22_X1 U2 ( .A1(n20), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U3 ( .A(b[31]), .ZN(n20) );
  INV_X1 U4 ( .A(n116), .ZN(n10) );
  INV_X1 U5 ( .A(n106), .ZN(n21) );
  INV_X1 U6 ( .A(n96), .ZN(n32) );
  AOI22_X1 U7 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U8 ( .A(n97), .ZN(n31) );
  INV_X1 U9 ( .A(n110), .ZN(n16) );
  INV_X1 U10 ( .A(n111), .ZN(n15) );
  INV_X1 U11 ( .A(n101), .ZN(n27) );
  INV_X1 U12 ( .A(n99), .ZN(n29) );
  INV_X1 U13 ( .A(n103), .ZN(n25) );
  INV_X1 U14 ( .A(n122), .ZN(n4) );
  INV_X1 U15 ( .A(n120), .ZN(n6) );
  INV_X1 U16 ( .A(n98), .ZN(n30) );
  AOI22_X1 U17 ( .A1(b[13]), .A2(a[13]), .B1(n19), .B2(n129), .ZN(n108) );
  INV_X1 U18 ( .A(n105), .ZN(n22) );
  INV_X1 U19 ( .A(n157), .ZN(n24) );
  AOI22_X1 U20 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n132), .ZN(n111) );
  INV_X1 U21 ( .A(n124), .ZN(n2) );
  AOI22_X1 U22 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  AOI22_X1 U23 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U24 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  INV_X1 U25 ( .A(n108), .ZN(n18) );
  AOI22_X1 U26 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  AOI22_X1 U27 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  AOI22_X1 U28 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  AOI22_X1 U29 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  INV_X1 U30 ( .A(n121), .ZN(n5) );
  AOI22_X1 U31 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  INV_X1 U32 ( .A(n123), .ZN(n3) );
  INV_X1 U33 ( .A(n118), .ZN(n8) );
  AOI22_X1 U34 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U35 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  INV_X1 U36 ( .A(n115), .ZN(n11) );
  INV_X1 U37 ( .A(n114), .ZN(n12) );
  INV_X1 U38 ( .A(n109), .ZN(n17) );
  INV_X1 U39 ( .A(n104), .ZN(n23) );
  INV_X1 U40 ( .A(n102), .ZN(n26) );
  INV_X1 U41 ( .A(n100), .ZN(n28) );
  AOI22_X1 U42 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U43 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  AOI22_X1 U44 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U45 ( .A1(b[15]), .A2(a[15]), .B1(n17), .B2(n131), .ZN(n110) );
  AOI22_X1 U46 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U47 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U48 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U49 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U50 ( .A1(b[14]), .A2(a[14]), .B1(n18), .B2(n130), .ZN(n109) );
  AOI22_X1 U51 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  AOI22_X1 U52 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  INV_X1 U53 ( .A(n119), .ZN(n7) );
  INV_X1 U54 ( .A(n117), .ZN(n9) );
  INV_X1 U55 ( .A(n113), .ZN(n13) );
  INV_X1 U56 ( .A(n112), .ZN(n14) );
  INV_X1 U57 ( .A(n107), .ZN(n19) );
  AOI22_X1 U58 ( .A1(b[12]), .A2(a[12]), .B1(n21), .B2(n128), .ZN(n107) );
  AOI22_X1 U59 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  AOI22_X1 U60 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  AOI22_X1 U61 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U62 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U63 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  XNOR2_X1 U64 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U65 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
endmodule


module carryLookAheadAdder_9 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n17), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n18), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n19), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n20), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n22), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n23), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  AOI22_X1 U1 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  INV_X1 U2 ( .A(a[31]), .ZN(n1) );
  OAI22_X1 U3 ( .A1(n21), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U4 ( .A(b[31]), .ZN(n21) );
  INV_X1 U5 ( .A(n117), .ZN(n9) );
  INV_X1 U6 ( .A(n108), .ZN(n18) );
  INV_X1 U7 ( .A(n96), .ZN(n32) );
  AOI22_X1 U8 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U9 ( .A(n110), .ZN(n16) );
  INV_X1 U10 ( .A(n97), .ZN(n31) );
  INV_X1 U11 ( .A(n103), .ZN(n25) );
  INV_X1 U12 ( .A(n109), .ZN(n17) );
  INV_X1 U13 ( .A(n106), .ZN(n20) );
  INV_X1 U14 ( .A(n102), .ZN(n26) );
  AOI22_X1 U15 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  INV_X1 U16 ( .A(n124), .ZN(n2) );
  AOI22_X1 U17 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  INV_X1 U18 ( .A(n112), .ZN(n14) );
  INV_X1 U19 ( .A(n113), .ZN(n13) );
  INV_X1 U20 ( .A(n99), .ZN(n29) );
  INV_X1 U21 ( .A(n100), .ZN(n28) );
  INV_X1 U22 ( .A(n122), .ZN(n4) );
  INV_X1 U23 ( .A(n119), .ZN(n7) );
  AOI22_X1 U24 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  INV_X1 U25 ( .A(n104), .ZN(n23) );
  INV_X1 U26 ( .A(n157), .ZN(n24) );
  AOI22_X1 U27 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  AOI22_X1 U28 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  INV_X1 U29 ( .A(n123), .ZN(n3) );
  XNOR2_X1 U30 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U31 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
  AOI22_X1 U32 ( .A1(b[15]), .A2(a[15]), .B1(n17), .B2(n131), .ZN(n110) );
  AOI22_X1 U33 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  AOI22_X1 U34 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  INV_X1 U35 ( .A(n107), .ZN(n19) );
  INV_X1 U36 ( .A(n101), .ZN(n27) );
  INV_X1 U37 ( .A(n121), .ZN(n5) );
  AOI22_X1 U38 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  AOI22_X1 U39 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  INV_X1 U40 ( .A(n118), .ZN(n8) );
  AOI22_X1 U41 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  INV_X1 U42 ( .A(n116), .ZN(n10) );
  AOI22_X1 U43 ( .A1(b[14]), .A2(a[14]), .B1(n18), .B2(n130), .ZN(n109) );
  AOI22_X1 U44 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  INV_X1 U45 ( .A(n111), .ZN(n15) );
  AOI22_X1 U46 ( .A1(b[11]), .A2(a[11]), .B1(n22), .B2(n127), .ZN(n106) );
  INV_X1 U47 ( .A(n98), .ZN(n30) );
  AOI22_X1 U48 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U49 ( .A1(b[12]), .A2(a[12]), .B1(n20), .B2(n128), .ZN(n107) );
  AOI22_X1 U50 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  AOI22_X1 U51 ( .A1(b[13]), .A2(a[13]), .B1(n19), .B2(n129), .ZN(n108) );
  AOI22_X1 U52 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U53 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U54 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U55 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  AOI22_X1 U56 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U57 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  AOI22_X1 U58 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  AOI22_X1 U59 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n132), .ZN(n111) );
  INV_X1 U60 ( .A(n120), .ZN(n6) );
  INV_X1 U61 ( .A(n115), .ZN(n11) );
  AOI22_X1 U62 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  INV_X1 U63 ( .A(n114), .ZN(n12) );
  INV_X1 U64 ( .A(n105), .ZN(n22) );
  AOI22_X1 U65 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
endmodule


module carryLookAheadAdder_8 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n26), .B(n155), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n28), .B(n153), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n30), .B(n151), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n17), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n18), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n19), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n20), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n21), .Z(result[11]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  INV_X1 U1 ( .A(n123), .ZN(n3) );
  AOI22_X1 U2 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  INV_X1 U3 ( .A(a[31]), .ZN(n1) );
  OAI22_X1 U4 ( .A1(n22), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U5 ( .A(b[31]), .ZN(n22) );
  INV_X1 U6 ( .A(n114), .ZN(n12) );
  INV_X1 U7 ( .A(n120), .ZN(n6) );
  AOI22_X1 U8 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  AOI22_X1 U9 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  XNOR2_X1 U10 ( .A(n104), .B(n126), .ZN(result[10]) );
  INV_X1 U11 ( .A(n99), .ZN(n29) );
  INV_X1 U12 ( .A(n108), .ZN(n18) );
  INV_X1 U13 ( .A(n110), .ZN(n16) );
  INV_X1 U14 ( .A(n103), .ZN(n25) );
  INV_X1 U15 ( .A(n106), .ZN(n20) );
  INV_X1 U16 ( .A(n96), .ZN(n32) );
  INV_X1 U17 ( .A(n97), .ZN(n31) );
  INV_X1 U18 ( .A(n112), .ZN(n14) );
  INV_X1 U19 ( .A(n101), .ZN(n27) );
  INV_X1 U20 ( .A(n102), .ZN(n26) );
  INV_X1 U21 ( .A(n105), .ZN(n21) );
  INV_X1 U22 ( .A(n98), .ZN(n30) );
  INV_X1 U23 ( .A(n122), .ZN(n4) );
  INV_X1 U24 ( .A(n118), .ZN(n8) );
  INV_X1 U25 ( .A(n116), .ZN(n10) );
  AOI22_X1 U26 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U27 ( .A1(b[13]), .A2(a[13]), .B1(n19), .B2(n129), .ZN(n108) );
  AOI22_X1 U28 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U29 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  INV_X1 U30 ( .A(n100), .ZN(n28) );
  AOI22_X1 U31 ( .A1(b[15]), .A2(a[15]), .B1(n17), .B2(n131), .ZN(n110) );
  AOI22_X1 U32 ( .A1(b[10]), .A2(a[10]), .B1(n23), .B2(n126), .ZN(n105) );
  AOI22_X1 U33 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U34 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  AOI22_X1 U35 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U36 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  AOI22_X1 U37 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  INV_X1 U38 ( .A(n121), .ZN(n5) );
  AOI22_X1 U39 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  AOI22_X1 U40 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U41 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U42 ( .A1(b[14]), .A2(a[14]), .B1(n18), .B2(n130), .ZN(n109) );
  AOI22_X1 U43 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U44 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  INV_X1 U45 ( .A(n111), .ZN(n15) );
  AOI22_X1 U46 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n132), .ZN(n111) );
  AOI22_X1 U47 ( .A1(b[11]), .A2(a[11]), .B1(n21), .B2(n127), .ZN(n106) );
  AOI22_X1 U48 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  AOI22_X1 U49 ( .A1(b[12]), .A2(a[12]), .B1(n20), .B2(n128), .ZN(n107) );
  AOI22_X1 U50 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U51 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  AOI22_X1 U52 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  INV_X1 U53 ( .A(n124), .ZN(n2) );
  AOI22_X1 U54 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  AOI22_X1 U55 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  INV_X1 U56 ( .A(n119), .ZN(n7) );
  INV_X1 U57 ( .A(n117), .ZN(n9) );
  INV_X1 U58 ( .A(n115), .ZN(n11) );
  INV_X1 U59 ( .A(n113), .ZN(n13) );
  INV_X1 U60 ( .A(n109), .ZN(n17) );
  INV_X1 U61 ( .A(n107), .ZN(n19) );
  INV_X1 U62 ( .A(n104), .ZN(n23) );
  INV_X1 U63 ( .A(n157), .ZN(n24) );
  AOI22_X1 U64 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  XNOR2_X1 U65 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U95 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
endmodule


module carryLookAheadAdder_7 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n17), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n18), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n19), .Z(result[13]) );
  XOR2_X1 U94 ( .A(n127), .B(n21), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n22), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  XOR2_X1 U1 ( .A(a[7]), .B(b[7]), .Z(n155) );
  INV_X1 U2 ( .A(a[31]), .ZN(n1) );
  OAI22_X1 U3 ( .A1(n23), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U4 ( .A(b[31]), .ZN(n23) );
  INV_X1 U5 ( .A(n119), .ZN(n7) );
  INV_X1 U6 ( .A(n108), .ZN(n18) );
  INV_X1 U7 ( .A(n124), .ZN(n2) );
  INV_X1 U8 ( .A(n104), .ZN(n22) );
  INV_X1 U9 ( .A(n122), .ZN(n4) );
  AOI22_X1 U10 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  INV_X1 U11 ( .A(n96), .ZN(n32) );
  XNOR2_X1 U12 ( .A(n106), .B(n128), .ZN(result[12]) );
  INV_X1 U13 ( .A(n97), .ZN(n31) );
  INV_X1 U14 ( .A(n98), .ZN(n30) );
  INV_X1 U15 ( .A(n99), .ZN(n29) );
  INV_X1 U16 ( .A(n103), .ZN(n25) );
  INV_X1 U17 ( .A(n113), .ZN(n13) );
  INV_X1 U18 ( .A(n109), .ZN(n17) );
  INV_X1 U19 ( .A(n112), .ZN(n14) );
  INV_X1 U20 ( .A(n107), .ZN(n19) );
  AOI22_X1 U21 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  INV_X1 U22 ( .A(n100), .ZN(n28) );
  AOI22_X1 U23 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  INV_X1 U24 ( .A(n105), .ZN(n21) );
  AOI22_X1 U25 ( .A1(b[15]), .A2(a[15]), .B1(n17), .B2(n131), .ZN(n110) );
  AOI22_X1 U26 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  AOI22_X1 U27 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U28 ( .A1(b[14]), .A2(a[14]), .B1(n18), .B2(n130), .ZN(n109) );
  AOI22_X1 U29 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U30 ( .A1(b[13]), .A2(a[13]), .B1(n19), .B2(n129), .ZN(n108) );
  INV_X1 U31 ( .A(n123), .ZN(n3) );
  AOI22_X1 U32 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  INV_X1 U33 ( .A(n115), .ZN(n11) );
  AOI22_X1 U34 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U35 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U36 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  INV_X1 U37 ( .A(n118), .ZN(n8) );
  INV_X1 U38 ( .A(n117), .ZN(n9) );
  INV_X1 U39 ( .A(n114), .ZN(n12) );
  AOI22_X1 U40 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  AOI22_X1 U41 ( .A1(b[10]), .A2(a[10]), .B1(n22), .B2(n126), .ZN(n105) );
  AOI22_X1 U42 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  AOI22_X1 U43 ( .A1(b[11]), .A2(a[11]), .B1(n21), .B2(n127), .ZN(n106) );
  AOI22_X1 U44 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U45 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  AOI22_X1 U46 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  AOI22_X1 U47 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  AOI22_X1 U48 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  AOI22_X1 U49 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  INV_X1 U50 ( .A(n121), .ZN(n5) );
  AOI22_X1 U51 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  INV_X1 U52 ( .A(n111), .ZN(n15) );
  AOI22_X1 U53 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  INV_X1 U54 ( .A(n102), .ZN(n26) );
  AOI22_X1 U55 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  INV_X1 U56 ( .A(n120), .ZN(n6) );
  AOI22_X1 U57 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  INV_X1 U58 ( .A(n116), .ZN(n10) );
  AOI22_X1 U59 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n132), .ZN(n111) );
  INV_X1 U60 ( .A(n110), .ZN(n16) );
  AOI22_X1 U61 ( .A1(b[12]), .A2(a[12]), .B1(n20), .B2(n128), .ZN(n107) );
  INV_X1 U62 ( .A(n106), .ZN(n20) );
  AOI22_X1 U63 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  INV_X1 U64 ( .A(n101), .ZN(n27) );
  INV_X1 U65 ( .A(n157), .ZN(n24) );
  XNOR2_X1 U93 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U121 ( .A1(b[9]), .A2(a[9]), .B1(n24), .B2(n158), .ZN(n104) );
endmodule


module carryLookAheadAdder_6 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n25), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n17), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n18), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n19), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n20), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n21), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n22), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  INV_X1 U1 ( .A(a[31]), .ZN(n1) );
  OAI22_X1 U2 ( .A1(n24), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U3 ( .A(b[31]), .ZN(n24) );
  INV_X1 U4 ( .A(n113), .ZN(n13) );
  INV_X1 U5 ( .A(n111), .ZN(n15) );
  INV_X1 U6 ( .A(n121), .ZN(n5) );
  INV_X1 U7 ( .A(n124), .ZN(n2) );
  INV_X1 U8 ( .A(n104), .ZN(n22) );
  AOI22_X1 U9 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  XNOR2_X1 U10 ( .A(n101), .B(n154), .ZN(result[6]) );
  INV_X1 U11 ( .A(n102), .ZN(n26) );
  INV_X1 U12 ( .A(n106), .ZN(n20) );
  INV_X1 U13 ( .A(n97), .ZN(n31) );
  AOI22_X1 U14 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  INV_X1 U15 ( .A(n96), .ZN(n32) );
  INV_X1 U16 ( .A(n105), .ZN(n21) );
  INV_X1 U17 ( .A(n98), .ZN(n30) );
  INV_X1 U18 ( .A(n100), .ZN(n28) );
  AOI22_X1 U19 ( .A1(b[11]), .A2(a[11]), .B1(n21), .B2(n127), .ZN(n106) );
  INV_X1 U20 ( .A(n107), .ZN(n19) );
  AOI22_X1 U21 ( .A1(b[10]), .A2(a[10]), .B1(n22), .B2(n126), .ZN(n105) );
  INV_X1 U22 ( .A(n115), .ZN(n11) );
  INV_X1 U23 ( .A(n122), .ZN(n4) );
  INV_X1 U24 ( .A(n119), .ZN(n7) );
  INV_X1 U25 ( .A(n116), .ZN(n10) );
  INV_X1 U26 ( .A(n109), .ZN(n17) );
  AOI22_X1 U27 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  INV_X1 U28 ( .A(n117), .ZN(n9) );
  AOI22_X1 U29 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U30 ( .A1(b[12]), .A2(a[12]), .B1(n20), .B2(n128), .ZN(n107) );
  AOI22_X1 U31 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U32 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  AOI22_X1 U33 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  AOI22_X1 U34 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  AOI22_X1 U35 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U36 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U37 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U38 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  AOI22_X1 U39 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U40 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  AOI22_X1 U41 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  AOI22_X1 U42 ( .A1(b[15]), .A2(a[15]), .B1(n17), .B2(n131), .ZN(n110) );
  AOI22_X1 U43 ( .A1(b[13]), .A2(a[13]), .B1(n19), .B2(n129), .ZN(n108) );
  AOI22_X1 U44 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  INV_X1 U45 ( .A(n123), .ZN(n3) );
  AOI22_X1 U46 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  INV_X1 U47 ( .A(n118), .ZN(n8) );
  AOI22_X1 U48 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  INV_X1 U49 ( .A(n120), .ZN(n6) );
  AOI22_X1 U50 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  INV_X1 U51 ( .A(n112), .ZN(n14) );
  AOI22_X1 U52 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  INV_X1 U53 ( .A(n114), .ZN(n12) );
  AOI22_X1 U54 ( .A1(b[14]), .A2(a[14]), .B1(n18), .B2(n130), .ZN(n109) );
  INV_X1 U55 ( .A(n108), .ZN(n18) );
  AOI22_X1 U56 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n132), .ZN(n111) );
  INV_X1 U57 ( .A(n110), .ZN(n16) );
  AOI22_X1 U58 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  INV_X1 U59 ( .A(n99), .ZN(n29) );
  AOI22_X1 U60 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  INV_X1 U61 ( .A(n101), .ZN(n27) );
  AOI22_X1 U62 ( .A1(b[8]), .A2(a[8]), .B1(n25), .B2(n156), .ZN(n157) );
  INV_X1 U63 ( .A(n103), .ZN(n25) );
  INV_X1 U64 ( .A(n157), .ZN(n23) );
  XNOR2_X1 U65 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U68 ( .A1(b[9]), .A2(a[9]), .B1(n23), .B2(n158), .ZN(n104) );
endmodule


module carryLookAheadAdder_5 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n24), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n26), .Z(result[7]) );
  XOR2_X1 U69 ( .A(n28), .B(n153), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n17), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n18), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n19), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n20), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n21), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n22), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  AOI22_X1 U1 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  INV_X1 U2 ( .A(a[31]), .ZN(n1) );
  OAI22_X1 U3 ( .A1(n25), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U4 ( .A(b[31]), .ZN(n25) );
  INV_X1 U5 ( .A(n115), .ZN(n11) );
  INV_X1 U6 ( .A(n110), .ZN(n16) );
  INV_X1 U7 ( .A(n124), .ZN(n2) );
  INV_X1 U8 ( .A(n120), .ZN(n6) );
  INV_X1 U9 ( .A(n96), .ZN(n32) );
  AOI22_X1 U10 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  XNOR2_X1 U11 ( .A(n101), .B(n154), .ZN(result[6]) );
  INV_X1 U12 ( .A(n106), .ZN(n20) );
  INV_X1 U13 ( .A(n112), .ZN(n14) );
  INV_X1 U14 ( .A(n104), .ZN(n22) );
  INV_X1 U15 ( .A(n97), .ZN(n31) );
  INV_X1 U16 ( .A(n116), .ZN(n10) );
  INV_X1 U17 ( .A(n100), .ZN(n28) );
  AOI22_X1 U18 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  INV_X1 U19 ( .A(n103), .ZN(n24) );
  INV_X1 U20 ( .A(n102), .ZN(n26) );
  INV_X1 U21 ( .A(n98), .ZN(n30) );
  AOI22_X1 U22 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  INV_X1 U23 ( .A(n157), .ZN(n23) );
  AOI22_X1 U24 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U25 ( .A1(b[7]), .A2(a[7]), .B1(n26), .B2(n155), .ZN(n103) );
  AOI22_X1 U26 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  AOI22_X1 U27 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U28 ( .A1(b[13]), .A2(a[13]), .B1(n19), .B2(n129), .ZN(n108) );
  AOI22_X1 U29 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  INV_X1 U30 ( .A(n101), .ZN(n27) );
  AOI22_X1 U31 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U32 ( .A1(b[14]), .A2(a[14]), .B1(n18), .B2(n130), .ZN(n109) );
  AOI22_X1 U33 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n132), .ZN(n111) );
  INV_X1 U34 ( .A(n119), .ZN(n7) );
  AOI22_X1 U35 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  INV_X1 U36 ( .A(n108), .ZN(n18) );
  INV_X1 U37 ( .A(n107), .ZN(n19) );
  INV_X1 U38 ( .A(n99), .ZN(n29) );
  AOI22_X1 U39 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U40 ( .A1(b[15]), .A2(a[15]), .B1(n17), .B2(n131), .ZN(n110) );
  AOI22_X1 U41 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  AOI22_X1 U42 ( .A1(b[8]), .A2(a[8]), .B1(n24), .B2(n156), .ZN(n157) );
  AOI22_X1 U43 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  AOI22_X1 U44 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  INV_X1 U45 ( .A(n105), .ZN(n21) );
  AOI22_X1 U46 ( .A1(b[10]), .A2(a[10]), .B1(n22), .B2(n126), .ZN(n105) );
  AOI22_X1 U47 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U48 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U49 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U50 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  INV_X1 U51 ( .A(n123), .ZN(n3) );
  INV_X1 U52 ( .A(n121), .ZN(n5) );
  INV_X1 U53 ( .A(n118), .ZN(n8) );
  INV_X1 U54 ( .A(n117), .ZN(n9) );
  INV_X1 U55 ( .A(n111), .ZN(n15) );
  AOI22_X1 U56 ( .A1(b[12]), .A2(a[12]), .B1(n20), .B2(n128), .ZN(n107) );
  INV_X1 U57 ( .A(n114), .ZN(n12) );
  INV_X1 U58 ( .A(n113), .ZN(n13) );
  INV_X1 U59 ( .A(n109), .ZN(n17) );
  AOI22_X1 U60 ( .A1(b[11]), .A2(a[11]), .B1(n21), .B2(n127), .ZN(n106) );
  AOI22_X1 U61 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  INV_X1 U62 ( .A(n122), .ZN(n4) );
  AOI22_X1 U63 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U64 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  XNOR2_X1 U65 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U68 ( .A1(b[9]), .A2(a[9]), .B1(n23), .B2(n158), .ZN(n104) );
endmodule


module carryLookAheadAdder_4 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n24), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n25), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n27), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n28), .Z(result[5]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n17), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n18), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n19), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n20), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n21), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n22), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  AOI22_X1 U1 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  INV_X1 U2 ( .A(n124), .ZN(n2) );
  INV_X1 U3 ( .A(a[31]), .ZN(n1) );
  OAI22_X1 U4 ( .A1(n26), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U5 ( .A(b[31]), .ZN(n26) );
  INV_X1 U6 ( .A(n122), .ZN(n4) );
  AOI22_X1 U7 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  INV_X1 U8 ( .A(n113), .ZN(n13) );
  INV_X1 U9 ( .A(n118), .ZN(n8) );
  INV_X1 U10 ( .A(n117), .ZN(n9) );
  INV_X1 U11 ( .A(n100), .ZN(n28) );
  INV_X1 U12 ( .A(n116), .ZN(n10) );
  INV_X1 U13 ( .A(n123), .ZN(n3) );
  AOI22_X1 U14 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  INV_X1 U15 ( .A(n96), .ZN(n32) );
  AOI22_X1 U16 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  AOI22_X1 U17 ( .A1(b[14]), .A2(a[14]), .B1(n18), .B2(n130), .ZN(n109) );
  XNOR2_X1 U18 ( .A(n99), .B(n152), .ZN(result[4]) );
  INV_X1 U19 ( .A(n103), .ZN(n24) );
  AOI22_X1 U20 ( .A1(b[8]), .A2(a[8]), .B1(n24), .B2(n156), .ZN(n157) );
  INV_X1 U21 ( .A(n109), .ZN(n17) );
  INV_X1 U22 ( .A(n112), .ZN(n14) );
  INV_X1 U23 ( .A(n108), .ZN(n18) );
  INV_X1 U24 ( .A(n97), .ZN(n31) );
  INV_X1 U25 ( .A(n98), .ZN(n30) );
  AOI22_X1 U26 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  INV_X1 U27 ( .A(n106), .ZN(n20) );
  INV_X1 U28 ( .A(n105), .ZN(n21) );
  INV_X1 U29 ( .A(n99), .ZN(n29) );
  AOI22_X1 U30 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U31 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  AOI22_X1 U32 ( .A1(b[15]), .A2(a[15]), .B1(n17), .B2(n131), .ZN(n110) );
  AOI22_X1 U33 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  INV_X1 U34 ( .A(n107), .ZN(n19) );
  AOI22_X1 U35 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U36 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  INV_X1 U37 ( .A(n119), .ZN(n7) );
  AOI22_X1 U38 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  AOI22_X1 U39 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U40 ( .A1(b[11]), .A2(a[11]), .B1(n21), .B2(n127), .ZN(n106) );
  AOI22_X1 U41 ( .A1(b[7]), .A2(a[7]), .B1(n25), .B2(n155), .ZN(n103) );
  AOI22_X1 U42 ( .A1(b[13]), .A2(a[13]), .B1(n19), .B2(n129), .ZN(n108) );
  AOI22_X1 U43 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U44 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  AOI22_X1 U45 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  AOI22_X1 U46 ( .A1(b[12]), .A2(a[12]), .B1(n20), .B2(n128), .ZN(n107) );
  AOI22_X1 U47 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U48 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  INV_X1 U49 ( .A(n121), .ZN(n5) );
  AOI22_X1 U50 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  INV_X1 U51 ( .A(n111), .ZN(n15) );
  AOI22_X1 U52 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n132), .ZN(n111) );
  INV_X1 U53 ( .A(n102), .ZN(n25) );
  AOI22_X1 U54 ( .A1(b[6]), .A2(a[6]), .B1(n27), .B2(n154), .ZN(n102) );
  AOI22_X1 U55 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  INV_X1 U56 ( .A(n115), .ZN(n11) );
  INV_X1 U57 ( .A(n120), .ZN(n6) );
  AOI22_X1 U58 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  INV_X1 U59 ( .A(n114), .ZN(n12) );
  INV_X1 U60 ( .A(n110), .ZN(n16) );
  AOI22_X1 U61 ( .A1(b[10]), .A2(a[10]), .B1(n22), .B2(n126), .ZN(n105) );
  INV_X1 U62 ( .A(n104), .ZN(n22) );
  INV_X1 U63 ( .A(n101), .ZN(n27) );
  INV_X1 U64 ( .A(n157), .ZN(n23) );
  XNOR2_X1 U65 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U70 ( .A1(b[9]), .A2(a[9]), .B1(n23), .B2(n158), .ZN(n104) );
endmodule


module carryLookAheadAdder_3 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n24), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n25), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n26), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n28), .B(n153), .Z(result[5]) );
  XOR2_X1 U71 ( .A(n30), .B(n151), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n17), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n18), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n19), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n20), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n21), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n22), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  XOR2_X1 U1 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U2 ( .A(a[3]), .B(b[3]), .Z(n151) );
  INV_X1 U3 ( .A(n108), .ZN(n18) );
  INV_X1 U4 ( .A(a[31]), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n27), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U6 ( .A(b[31]), .ZN(n27) );
  INV_X1 U7 ( .A(n107), .ZN(n19) );
  INV_X1 U8 ( .A(n114), .ZN(n12) );
  INV_X1 U9 ( .A(n116), .ZN(n10) );
  INV_X1 U10 ( .A(n120), .ZN(n6) );
  INV_X1 U11 ( .A(n96), .ZN(n32) );
  AOI22_X1 U12 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  XNOR2_X1 U13 ( .A(n99), .B(n152), .ZN(result[4]) );
  INV_X1 U14 ( .A(n99), .ZN(n29) );
  INV_X1 U15 ( .A(n97), .ZN(n31) );
  INV_X1 U16 ( .A(n98), .ZN(n30) );
  INV_X1 U17 ( .A(n106), .ZN(n20) );
  INV_X1 U18 ( .A(n101), .ZN(n26) );
  INV_X1 U19 ( .A(n102), .ZN(n25) );
  INV_X1 U20 ( .A(n103), .ZN(n24) );
  AOI22_X1 U21 ( .A1(b[8]), .A2(a[8]), .B1(n24), .B2(n156), .ZN(n157) );
  AOI22_X1 U22 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U23 ( .A1(b[7]), .A2(a[7]), .B1(n25), .B2(n155), .ZN(n103) );
  AOI22_X1 U24 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  AOI22_X1 U25 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  AOI22_X1 U26 ( .A1(b[5]), .A2(a[5]), .B1(n28), .B2(n153), .ZN(n101) );
  AOI22_X1 U27 ( .A1(b[15]), .A2(a[15]), .B1(n17), .B2(n131), .ZN(n110) );
  AOI22_X1 U28 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  INV_X1 U29 ( .A(n118), .ZN(n8) );
  AOI22_X1 U30 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  INV_X1 U31 ( .A(n123), .ZN(n3) );
  AOI22_X1 U32 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U33 ( .A1(b[10]), .A2(a[10]), .B1(n22), .B2(n126), .ZN(n105) );
  INV_X1 U34 ( .A(n113), .ZN(n13) );
  AOI22_X1 U35 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  AOI22_X1 U36 ( .A1(b[13]), .A2(a[13]), .B1(n19), .B2(n129), .ZN(n108) );
  INV_X1 U37 ( .A(n124), .ZN(n2) );
  AOI22_X1 U38 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  AOI22_X1 U39 ( .A1(b[6]), .A2(a[6]), .B1(n26), .B2(n154), .ZN(n102) );
  AOI22_X1 U40 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  INV_X1 U41 ( .A(n112), .ZN(n14) );
  INV_X1 U42 ( .A(n110), .ZN(n16) );
  AOI22_X1 U43 ( .A1(b[14]), .A2(a[14]), .B1(n18), .B2(n130), .ZN(n109) );
  AOI22_X1 U44 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  AOI22_X1 U45 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U46 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U47 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  AOI22_X1 U48 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n132), .ZN(n111) );
  AOI22_X1 U49 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  AOI22_X1 U50 ( .A1(b[12]), .A2(a[12]), .B1(n20), .B2(n128), .ZN(n107) );
  AOI22_X1 U51 ( .A1(b[11]), .A2(a[11]), .B1(n21), .B2(n127), .ZN(n106) );
  AOI22_X1 U52 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U53 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  AOI22_X1 U54 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  INV_X1 U55 ( .A(n122), .ZN(n4) );
  INV_X1 U56 ( .A(n121), .ZN(n5) );
  INV_X1 U57 ( .A(n119), .ZN(n7) );
  INV_X1 U58 ( .A(n117), .ZN(n9) );
  INV_X1 U59 ( .A(n115), .ZN(n11) );
  INV_X1 U60 ( .A(n111), .ZN(n15) );
  INV_X1 U61 ( .A(n109), .ZN(n17) );
  INV_X1 U62 ( .A(n105), .ZN(n21) );
  INV_X1 U63 ( .A(n104), .ZN(n22) );
  INV_X1 U64 ( .A(n157), .ZN(n23) );
  INV_X1 U65 ( .A(n100), .ZN(n28) );
  AOI22_X1 U70 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  XNOR2_X1 U120 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U125 ( .A1(b[9]), .A2(a[9]), .B1(n23), .B2(n158), .ZN(n104) );
endmodule


module carryLookAheadAdder_2 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n24), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n25), .Z(result[7]) );
  XOR2_X1 U69 ( .A(n27), .B(n153), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n17), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n18), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n19), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n20), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n21), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n22), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  XOR2_X1 U1 ( .A(a[5]), .B(b[5]), .Z(n153) );
  INV_X1 U2 ( .A(n106), .ZN(n20) );
  AOI22_X1 U3 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  INV_X1 U4 ( .A(a[31]), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n28), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U6 ( .A(b[31]), .ZN(n28) );
  INV_X1 U7 ( .A(n118), .ZN(n8) );
  INV_X1 U8 ( .A(n120), .ZN(n6) );
  INV_X1 U9 ( .A(n114), .ZN(n12) );
  AOI22_X1 U10 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  XNOR2_X1 U11 ( .A(n101), .B(n154), .ZN(result[6]) );
  INV_X1 U12 ( .A(n101), .ZN(n26) );
  INV_X1 U13 ( .A(n96), .ZN(n32) );
  INV_X1 U14 ( .A(n97), .ZN(n31) );
  INV_X1 U15 ( .A(n99), .ZN(n29) );
  INV_X1 U16 ( .A(n108), .ZN(n18) );
  INV_X1 U17 ( .A(n157), .ZN(n23) );
  AOI22_X1 U18 ( .A1(b[8]), .A2(a[8]), .B1(n24), .B2(n156), .ZN(n157) );
  INV_X1 U19 ( .A(n107), .ZN(n19) );
  AOI22_X1 U20 ( .A1(b[5]), .A2(a[5]), .B1(n27), .B2(n153), .ZN(n101) );
  INV_X1 U21 ( .A(n123), .ZN(n3) );
  INV_X1 U22 ( .A(n103), .ZN(n24) );
  AOI22_X1 U23 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U24 ( .A1(b[15]), .A2(a[15]), .B1(n17), .B2(n131), .ZN(n110) );
  AOI22_X1 U25 ( .A1(b[13]), .A2(a[13]), .B1(n19), .B2(n129), .ZN(n108) );
  AOI22_X1 U26 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  AOI22_X1 U27 ( .A1(b[14]), .A2(a[14]), .B1(n18), .B2(n130), .ZN(n109) );
  INV_X1 U28 ( .A(n100), .ZN(n27) );
  AOI22_X1 U29 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  INV_X1 U30 ( .A(n110), .ZN(n16) );
  INV_X1 U31 ( .A(n98), .ZN(n30) );
  AOI22_X1 U32 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U33 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  AOI22_X1 U34 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U35 ( .A1(b[12]), .A2(a[12]), .B1(n20), .B2(n128), .ZN(n107) );
  AOI22_X1 U36 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  AOI22_X1 U37 ( .A1(b[6]), .A2(a[6]), .B1(n26), .B2(n154), .ZN(n102) );
  AOI22_X1 U38 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U39 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n132), .ZN(n111) );
  AOI22_X1 U40 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U41 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  AOI22_X1 U42 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  INV_X1 U43 ( .A(n122), .ZN(n4) );
  AOI22_X1 U44 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  INV_X1 U45 ( .A(n124), .ZN(n2) );
  AOI22_X1 U46 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  INV_X1 U47 ( .A(n119), .ZN(n7) );
  INV_X1 U48 ( .A(n117), .ZN(n9) );
  INV_X1 U49 ( .A(n113), .ZN(n13) );
  INV_X1 U50 ( .A(n112), .ZN(n14) );
  INV_X1 U51 ( .A(n109), .ZN(n17) );
  AOI22_X1 U52 ( .A1(b[11]), .A2(a[11]), .B1(n21), .B2(n127), .ZN(n106) );
  AOI22_X1 U53 ( .A1(b[10]), .A2(a[10]), .B1(n22), .B2(n126), .ZN(n105) );
  AOI22_X1 U54 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  AOI22_X1 U55 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  AOI22_X1 U56 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  INV_X1 U57 ( .A(n121), .ZN(n5) );
  INV_X1 U58 ( .A(n116), .ZN(n10) );
  INV_X1 U59 ( .A(n115), .ZN(n11) );
  AOI22_X1 U60 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  INV_X1 U61 ( .A(n111), .ZN(n15) );
  INV_X1 U62 ( .A(n105), .ZN(n21) );
  INV_X1 U63 ( .A(n104), .ZN(n22) );
  AOI22_X1 U64 ( .A1(b[7]), .A2(a[7]), .B1(n25), .B2(n155), .ZN(n103) );
  INV_X1 U65 ( .A(n102), .ZN(n25) );
  XNOR2_X1 U68 ( .A(n158), .B(n157), .ZN(result[9]) );
  AOI22_X1 U123 ( .A1(b[9]), .A2(a[9]), .B1(n23), .B2(n158), .ZN(n104) );
endmodule


module carryLookAheadAdder_1 ( a, b, cin, result, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  input cin;
  output cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158;

  XOR2_X1 U66 ( .A(n24), .B(n156), .Z(result[8]) );
  XOR2_X1 U67 ( .A(n155), .B(n25), .Z(result[7]) );
  XOR2_X1 U68 ( .A(n26), .B(n154), .Z(result[6]) );
  XOR2_X1 U69 ( .A(n153), .B(n27), .Z(result[5]) );
  XOR2_X1 U70 ( .A(n29), .B(n152), .Z(result[4]) );
  XOR2_X1 U71 ( .A(n151), .B(n30), .Z(result[3]) );
  XOR2_X1 U72 ( .A(n150), .B(n149), .Z(result[31]) );
  XOR2_X1 U73 ( .A(n2), .B(n148), .Z(result[30]) );
  XOR2_X1 U74 ( .A(n31), .B(n147), .Z(result[2]) );
  XOR2_X1 U75 ( .A(n146), .B(n3), .Z(result[29]) );
  XOR2_X1 U76 ( .A(n4), .B(n145), .Z(result[28]) );
  XOR2_X1 U77 ( .A(n144), .B(n5), .Z(result[27]) );
  XOR2_X1 U78 ( .A(n6), .B(n143), .Z(result[26]) );
  XOR2_X1 U79 ( .A(n142), .B(n7), .Z(result[25]) );
  XOR2_X1 U80 ( .A(n8), .B(n141), .Z(result[24]) );
  XOR2_X1 U81 ( .A(n140), .B(n9), .Z(result[23]) );
  XOR2_X1 U82 ( .A(n10), .B(n139), .Z(result[22]) );
  XOR2_X1 U83 ( .A(n138), .B(n11), .Z(result[21]) );
  XOR2_X1 U84 ( .A(n12), .B(n137), .Z(result[20]) );
  XOR2_X1 U85 ( .A(n136), .B(n32), .Z(result[1]) );
  XOR2_X1 U86 ( .A(n135), .B(n13), .Z(result[19]) );
  XOR2_X1 U87 ( .A(n14), .B(n134), .Z(result[18]) );
  XOR2_X1 U88 ( .A(n133), .B(n15), .Z(result[17]) );
  XOR2_X1 U89 ( .A(n16), .B(n132), .Z(result[16]) );
  XOR2_X1 U90 ( .A(n131), .B(n17), .Z(result[15]) );
  XOR2_X1 U91 ( .A(n18), .B(n130), .Z(result[14]) );
  XOR2_X1 U92 ( .A(n129), .B(n19), .Z(result[13]) );
  XOR2_X1 U93 ( .A(n20), .B(n128), .Z(result[12]) );
  XOR2_X1 U94 ( .A(n127), .B(n21), .Z(result[11]) );
  XOR2_X1 U95 ( .A(n22), .B(n126), .Z(result[10]) );
  XOR2_X1 U96 ( .A(cin), .B(n125), .Z(result[0]) );
  XOR2_X1 U97 ( .A(n1), .B(b[31]), .Z(n150) );
  XOR2_X1 U98 ( .A(a[30]), .B(b[30]), .Z(n148) );
  XOR2_X1 U99 ( .A(a[29]), .B(b[29]), .Z(n146) );
  XOR2_X1 U100 ( .A(a[28]), .B(b[28]), .Z(n145) );
  XOR2_X1 U101 ( .A(a[27]), .B(b[27]), .Z(n144) );
  XOR2_X1 U102 ( .A(a[26]), .B(b[26]), .Z(n143) );
  XOR2_X1 U103 ( .A(a[25]), .B(b[25]), .Z(n142) );
  XOR2_X1 U104 ( .A(a[24]), .B(b[24]), .Z(n141) );
  XOR2_X1 U105 ( .A(a[23]), .B(b[23]), .Z(n140) );
  XOR2_X1 U106 ( .A(a[22]), .B(b[22]), .Z(n139) );
  XOR2_X1 U107 ( .A(a[21]), .B(b[21]), .Z(n138) );
  XOR2_X1 U108 ( .A(a[20]), .B(b[20]), .Z(n137) );
  XOR2_X1 U109 ( .A(a[19]), .B(b[19]), .Z(n135) );
  XOR2_X1 U110 ( .A(a[18]), .B(b[18]), .Z(n134) );
  XOR2_X1 U111 ( .A(a[17]), .B(b[17]), .Z(n133) );
  XOR2_X1 U112 ( .A(a[16]), .B(b[16]), .Z(n132) );
  XOR2_X1 U113 ( .A(a[15]), .B(b[15]), .Z(n131) );
  XOR2_X1 U114 ( .A(a[14]), .B(b[14]), .Z(n130) );
  XOR2_X1 U115 ( .A(a[13]), .B(b[13]), .Z(n129) );
  XOR2_X1 U116 ( .A(a[12]), .B(b[12]), .Z(n128) );
  XOR2_X1 U117 ( .A(a[11]), .B(b[11]), .Z(n127) );
  XOR2_X1 U118 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U119 ( .A(a[9]), .B(b[9]), .Z(n158) );
  XOR2_X1 U120 ( .A(a[8]), .B(b[8]), .Z(n156) );
  XOR2_X1 U121 ( .A(a[7]), .B(b[7]), .Z(n155) );
  XOR2_X1 U122 ( .A(a[6]), .B(b[6]), .Z(n154) );
  XOR2_X1 U123 ( .A(a[5]), .B(b[5]), .Z(n153) );
  XOR2_X1 U124 ( .A(a[4]), .B(b[4]), .Z(n152) );
  XOR2_X1 U125 ( .A(a[3]), .B(b[3]), .Z(n151) );
  XOR2_X1 U126 ( .A(a[2]), .B(b[2]), .Z(n147) );
  XOR2_X1 U127 ( .A(a[1]), .B(b[1]), .Z(n136) );
  XOR2_X1 U128 ( .A(a[0]), .B(b[0]), .Z(n125) );
  AOI22_X1 U1 ( .A1(b[30]), .A2(a[30]), .B1(n2), .B2(n148), .ZN(n149) );
  INV_X1 U2 ( .A(a[31]), .ZN(n1) );
  INV_X1 U3 ( .A(n110), .ZN(n16) );
  INV_X1 U4 ( .A(n116), .ZN(n10) );
  INV_X1 U5 ( .A(n104), .ZN(n22) );
  OAI22_X1 U6 ( .A1(n28), .A2(n1), .B1(n149), .B2(n150), .ZN(cout) );
  INV_X1 U7 ( .A(b[31]), .ZN(n28) );
  INV_X1 U8 ( .A(n96), .ZN(n32) );
  INV_X1 U9 ( .A(n97), .ZN(n31) );
  INV_X1 U10 ( .A(n99), .ZN(n29) );
  AOI22_X1 U11 ( .A1(b[8]), .A2(a[8]), .B1(n24), .B2(n156), .ZN(n157) );
  INV_X1 U12 ( .A(n118), .ZN(n8) );
  AOI22_X1 U13 ( .A1(b[0]), .A2(a[0]), .B1(n125), .B2(cin), .ZN(n96) );
  AOI22_X1 U14 ( .A1(b[1]), .A2(a[1]), .B1(n32), .B2(n136), .ZN(n97) );
  AOI22_X1 U15 ( .A1(b[19]), .A2(a[19]), .B1(n13), .B2(n135), .ZN(n114) );
  AOI22_X1 U16 ( .A1(b[10]), .A2(a[10]), .B1(n22), .B2(n126), .ZN(n105) );
  INV_X1 U17 ( .A(n103), .ZN(n24) );
  AOI22_X1 U18 ( .A1(b[3]), .A2(a[3]), .B1(n30), .B2(n151), .ZN(n99) );
  AOI22_X1 U19 ( .A1(b[9]), .A2(a[9]), .B1(n23), .B2(n158), .ZN(n104) );
  AOI22_X1 U20 ( .A1(b[7]), .A2(a[7]), .B1(n25), .B2(n155), .ZN(n103) );
  AOI22_X1 U21 ( .A1(b[6]), .A2(a[6]), .B1(n26), .B2(n154), .ZN(n102) );
  AOI22_X1 U22 ( .A1(b[13]), .A2(a[13]), .B1(n19), .B2(n129), .ZN(n108) );
  INV_X1 U23 ( .A(n106), .ZN(n20) );
  INV_X1 U24 ( .A(n101), .ZN(n26) );
  AOI22_X1 U25 ( .A1(b[4]), .A2(a[4]), .B1(n29), .B2(n152), .ZN(n100) );
  AOI22_X1 U26 ( .A1(b[12]), .A2(a[12]), .B1(n20), .B2(n128), .ZN(n107) );
  AOI22_X1 U27 ( .A1(b[21]), .A2(a[21]), .B1(n11), .B2(n138), .ZN(n116) );
  AOI22_X1 U28 ( .A1(b[16]), .A2(a[16]), .B1(n16), .B2(n132), .ZN(n111) );
  AOI22_X1 U29 ( .A1(b[11]), .A2(a[11]), .B1(n21), .B2(n127), .ZN(n106) );
  AOI22_X1 U30 ( .A1(b[5]), .A2(a[5]), .B1(n27), .B2(n153), .ZN(n101) );
  AOI22_X1 U31 ( .A1(b[20]), .A2(a[20]), .B1(n12), .B2(n137), .ZN(n115) );
  AOI22_X1 U32 ( .A1(b[15]), .A2(a[15]), .B1(n17), .B2(n131), .ZN(n110) );
  XNOR2_X1 U33 ( .A(n158), .B(n157), .ZN(result[9]) );
  INV_X1 U34 ( .A(n157), .ZN(n23) );
  INV_X1 U35 ( .A(n102), .ZN(n25) );
  INV_X1 U36 ( .A(n100), .ZN(n27) );
  INV_X1 U37 ( .A(n98), .ZN(n30) );
  AOI22_X1 U38 ( .A1(b[2]), .A2(a[2]), .B1(n31), .B2(n147), .ZN(n98) );
  AOI22_X1 U39 ( .A1(b[18]), .A2(a[18]), .B1(n14), .B2(n134), .ZN(n113) );
  AOI22_X1 U40 ( .A1(b[17]), .A2(a[17]), .B1(n15), .B2(n133), .ZN(n112) );
  AOI22_X1 U41 ( .A1(b[23]), .A2(a[23]), .B1(n9), .B2(n140), .ZN(n118) );
  INV_X1 U42 ( .A(n112), .ZN(n14) );
  AOI22_X1 U43 ( .A1(b[14]), .A2(a[14]), .B1(n18), .B2(n130), .ZN(n109) );
  AOI22_X1 U44 ( .A1(b[25]), .A2(a[25]), .B1(n7), .B2(n142), .ZN(n120) );
  AOI22_X1 U45 ( .A1(b[26]), .A2(a[26]), .B1(n6), .B2(n143), .ZN(n121) );
  AOI22_X1 U46 ( .A1(b[27]), .A2(a[27]), .B1(n5), .B2(n144), .ZN(n122) );
  INV_X1 U47 ( .A(n119), .ZN(n7) );
  INV_X1 U48 ( .A(n114), .ZN(n12) );
  INV_X1 U49 ( .A(n109), .ZN(n17) );
  INV_X1 U50 ( .A(n108), .ZN(n18) );
  INV_X1 U51 ( .A(n120), .ZN(n6) );
  AOI22_X1 U52 ( .A1(b[24]), .A2(a[24]), .B1(n8), .B2(n141), .ZN(n119) );
  AOI22_X1 U53 ( .A1(b[22]), .A2(a[22]), .B1(n10), .B2(n139), .ZN(n117) );
  INV_X1 U54 ( .A(n122), .ZN(n4) );
  AOI22_X1 U55 ( .A1(b[28]), .A2(a[28]), .B1(n4), .B2(n145), .ZN(n123) );
  INV_X1 U56 ( .A(n124), .ZN(n2) );
  AOI22_X1 U57 ( .A1(b[29]), .A2(a[29]), .B1(n3), .B2(n146), .ZN(n124) );
  INV_X1 U58 ( .A(n123), .ZN(n3) );
  INV_X1 U59 ( .A(n121), .ZN(n5) );
  INV_X1 U60 ( .A(n117), .ZN(n9) );
  INV_X1 U61 ( .A(n115), .ZN(n11) );
  INV_X1 U62 ( .A(n113), .ZN(n13) );
  INV_X1 U63 ( .A(n111), .ZN(n15) );
  INV_X1 U64 ( .A(n107), .ZN(n19) );
  INV_X1 U65 ( .A(n105), .ZN(n21) );
endmodule


module multiplierTreeV2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n56, n58,
         n60, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n89, n90, n91, n92,
         n93, n94, n95, n100;
  wire   [63:1] carry;

  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .S(SUM[0]) );
  FA_X1 U1_62 ( .A(A[62]), .B(1'b0), .CI(n2), .CO(carry[63]), .S(SUM[62]) );
  XNOR2_X2 U1 ( .A(A[63]), .B(carry[63]), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(SUM[63]) );
  AND2_X1 U3 ( .A1(A[61]), .A2(n13), .ZN(n2) );
  AND2_X1 U4 ( .A1(A[52]), .A2(n5), .ZN(n3) );
  AND2_X1 U5 ( .A1(A[53]), .A2(n3), .ZN(n4) );
  AND2_X1 U6 ( .A1(A[51]), .A2(n7), .ZN(n5) );
  AND2_X1 U7 ( .A1(A[57]), .A2(n8), .ZN(n6) );
  AND2_X1 U8 ( .A1(A[50]), .A2(n14), .ZN(n7) );
  AND2_X1 U9 ( .A1(A[56]), .A2(n10), .ZN(n8) );
  AND2_X1 U10 ( .A1(A[58]), .A2(n6), .ZN(n9) );
  AND2_X1 U11 ( .A1(A[55]), .A2(n11), .ZN(n10) );
  AND2_X1 U12 ( .A1(A[54]), .A2(n4), .ZN(n11) );
  AND2_X1 U13 ( .A1(A[59]), .A2(n9), .ZN(n12) );
  AND2_X1 U14 ( .A1(A[60]), .A2(n12), .ZN(n13) );
  AND2_X1 U15 ( .A1(A[49]), .A2(n15), .ZN(n14) );
  AND2_X1 U16 ( .A1(A[48]), .A2(n21), .ZN(n15) );
  AND2_X1 U17 ( .A1(A[39]), .A2(n18), .ZN(n16) );
  AND2_X1 U18 ( .A1(A[36]), .A2(n19), .ZN(n17) );
  AND2_X1 U19 ( .A1(A[38]), .A2(n20), .ZN(n18) );
  AND2_X1 U20 ( .A1(A[35]), .A2(n56), .ZN(n19) );
  AND2_X1 U21 ( .A1(A[37]), .A2(n17), .ZN(n20) );
  AND2_X1 U22 ( .A1(A[47]), .A2(n26), .ZN(n21) );
  AND2_X1 U23 ( .A1(A[42]), .A2(n25), .ZN(n22) );
  AND2_X1 U24 ( .A1(A[43]), .A2(n22), .ZN(n23) );
  AND2_X1 U25 ( .A1(A[40]), .A2(n16), .ZN(n24) );
  AND2_X1 U26 ( .A1(A[41]), .A2(n24), .ZN(n25) );
  AND2_X1 U27 ( .A1(A[46]), .A2(n28), .ZN(n26) );
  AND2_X1 U28 ( .A1(A[44]), .A2(n23), .ZN(n27) );
  AND2_X1 U29 ( .A1(A[45]), .A2(n27), .ZN(n28) );
  XOR2_X1 U30 ( .A(A[57]), .B(n8), .Z(SUM[57]) );
  XOR2_X1 U31 ( .A(A[58]), .B(n6), .Z(SUM[58]) );
  XOR2_X1 U32 ( .A(A[59]), .B(n9), .Z(SUM[59]) );
  XOR2_X1 U33 ( .A(A[61]), .B(n13), .Z(SUM[61]) );
  XOR2_X1 U34 ( .A(A[60]), .B(n12), .Z(SUM[60]) );
  XOR2_X1 U35 ( .A(A[47]), .B(n26), .Z(SUM[47]) );
  XOR2_X1 U36 ( .A(A[48]), .B(n21), .Z(SUM[48]) );
  XOR2_X1 U37 ( .A(A[49]), .B(n15), .Z(SUM[49]) );
  XOR2_X1 U38 ( .A(A[50]), .B(n14), .Z(SUM[50]) );
  XOR2_X1 U39 ( .A(A[51]), .B(n7), .Z(SUM[51]) );
  XOR2_X1 U40 ( .A(A[52]), .B(n5), .Z(SUM[52]) );
  XOR2_X1 U41 ( .A(A[53]), .B(n3), .Z(SUM[53]) );
  XOR2_X1 U42 ( .A(A[54]), .B(n4), .Z(SUM[54]) );
  XOR2_X1 U43 ( .A(A[55]), .B(n11), .Z(SUM[55]) );
  XOR2_X1 U44 ( .A(A[56]), .B(n10), .Z(SUM[56]) );
  XOR2_X1 U45 ( .A(A[35]), .B(n56), .Z(SUM[35]) );
  XOR2_X1 U46 ( .A(A[36]), .B(n19), .Z(SUM[36]) );
  XOR2_X1 U47 ( .A(A[37]), .B(n17), .Z(SUM[37]) );
  XOR2_X1 U48 ( .A(A[38]), .B(n20), .Z(SUM[38]) );
  XOR2_X1 U49 ( .A(A[39]), .B(n18), .Z(SUM[39]) );
  XOR2_X1 U50 ( .A(A[40]), .B(n16), .Z(SUM[40]) );
  XOR2_X1 U51 ( .A(A[41]), .B(n24), .Z(SUM[41]) );
  XOR2_X1 U52 ( .A(A[42]), .B(n25), .Z(SUM[42]) );
  XOR2_X1 U53 ( .A(A[43]), .B(n22), .Z(SUM[43]) );
  XOR2_X1 U54 ( .A(A[44]), .B(n23), .Z(SUM[44]) );
  XOR2_X1 U55 ( .A(A[45]), .B(n27), .Z(SUM[45]) );
  XOR2_X1 U56 ( .A(A[46]), .B(n28), .Z(SUM[46]) );
  AND2_X1 U57 ( .A1(A[34]), .A2(n58), .ZN(n56) );
  XOR2_X1 U58 ( .A(A[34]), .B(n58), .Z(SUM[34]) );
  AND2_X1 U59 ( .A1(A[33]), .A2(n60), .ZN(n58) );
  XOR2_X1 U60 ( .A(A[33]), .B(n60), .Z(SUM[33]) );
  AND2_X1 U61 ( .A1(A[32]), .A2(n64), .ZN(n60) );
  XOR2_X1 U62 ( .A(A[32]), .B(n64), .Z(SUM[32]) );
  AND2_X1 U63 ( .A1(A[28]), .A2(n70), .ZN(n62) );
  AND2_X1 U64 ( .A1(A[29]), .A2(n62), .ZN(n63) );
  AND2_X1 U65 ( .A1(A[31]), .A2(n65), .ZN(n64) );
  AND2_X1 U66 ( .A1(A[30]), .A2(n63), .ZN(n65) );
  AND2_X1 U67 ( .A1(A[23]), .A2(n77), .ZN(n66) );
  AND2_X1 U68 ( .A1(A[24]), .A2(n66), .ZN(n67) );
  AND2_X1 U69 ( .A1(A[25]), .A2(n67), .ZN(n68) );
  AND2_X1 U70 ( .A1(A[26]), .A2(n68), .ZN(n69) );
  AND2_X1 U71 ( .A1(A[27]), .A2(n69), .ZN(n70) );
  AND2_X1 U72 ( .A1(A[16]), .A2(n84), .ZN(n71) );
  AND2_X1 U73 ( .A1(A[17]), .A2(n71), .ZN(n72) );
  AND2_X1 U74 ( .A1(A[18]), .A2(n72), .ZN(n73) );
  AND2_X1 U75 ( .A1(A[19]), .A2(n73), .ZN(n74) );
  AND2_X1 U76 ( .A1(A[20]), .A2(n74), .ZN(n75) );
  AND2_X1 U77 ( .A1(A[21]), .A2(n75), .ZN(n76) );
  AND2_X1 U78 ( .A1(A[22]), .A2(n76), .ZN(n77) );
  AND2_X1 U79 ( .A1(A[9]), .A2(n95), .ZN(n78) );
  AND2_X1 U80 ( .A1(A[10]), .A2(n78), .ZN(n79) );
  AND2_X1 U81 ( .A1(A[11]), .A2(n79), .ZN(n80) );
  AND2_X1 U82 ( .A1(A[12]), .A2(n80), .ZN(n81) );
  AND2_X1 U83 ( .A1(A[13]), .A2(n81), .ZN(n82) );
  AND2_X1 U84 ( .A1(A[14]), .A2(n82), .ZN(n83) );
  AND2_X1 U85 ( .A1(A[15]), .A2(n83), .ZN(n84) );
  XOR2_X1 U86 ( .A(A[28]), .B(n70), .Z(SUM[28]) );
  XOR2_X1 U87 ( .A(A[29]), .B(n62), .Z(SUM[29]) );
  XOR2_X1 U88 ( .A(A[30]), .B(n63), .Z(SUM[30]) );
  XOR2_X1 U89 ( .A(A[31]), .B(n65), .Z(SUM[31]) );
  AND2_X1 U90 ( .A1(A[2]), .A2(n100), .ZN(n89) );
  AND2_X1 U91 ( .A1(A[3]), .A2(n89), .ZN(n90) );
  AND2_X1 U92 ( .A1(A[4]), .A2(n90), .ZN(n91) );
  AND2_X1 U93 ( .A1(A[5]), .A2(n91), .ZN(n92) );
  AND2_X1 U94 ( .A1(A[6]), .A2(n92), .ZN(n93) );
  AND2_X1 U95 ( .A1(A[7]), .A2(n93), .ZN(n94) );
  AND2_X1 U96 ( .A1(A[8]), .A2(n94), .ZN(n95) );
  XOR2_X1 U97 ( .A(A[26]), .B(n68), .Z(SUM[26]) );
  XOR2_X1 U98 ( .A(A[27]), .B(n69), .Z(SUM[27]) );
  XOR2_X1 U99 ( .A(A[24]), .B(n66), .Z(SUM[24]) );
  XOR2_X1 U100 ( .A(A[25]), .B(n67), .Z(SUM[25]) );
  AND2_X1 U101 ( .A1(A[1]), .A2(carry[1]), .ZN(n100) );
  XOR2_X1 U102 ( .A(A[19]), .B(n73), .Z(SUM[19]) );
  XOR2_X1 U103 ( .A(A[20]), .B(n74), .Z(SUM[20]) );
  XOR2_X1 U104 ( .A(A[21]), .B(n75), .Z(SUM[21]) );
  XOR2_X1 U105 ( .A(A[22]), .B(n76), .Z(SUM[22]) );
  XOR2_X1 U106 ( .A(A[23]), .B(n77), .Z(SUM[23]) );
  XOR2_X1 U107 ( .A(A[15]), .B(n83), .Z(SUM[15]) );
  XOR2_X1 U108 ( .A(A[16]), .B(n84), .Z(SUM[16]) );
  XOR2_X1 U109 ( .A(A[17]), .B(n71), .Z(SUM[17]) );
  XOR2_X1 U110 ( .A(A[18]), .B(n72), .Z(SUM[18]) );
  XOR2_X1 U111 ( .A(A[11]), .B(n79), .Z(SUM[11]) );
  XOR2_X1 U112 ( .A(A[12]), .B(n80), .Z(SUM[12]) );
  XOR2_X1 U113 ( .A(A[13]), .B(n81), .Z(SUM[13]) );
  XOR2_X1 U114 ( .A(A[14]), .B(n82), .Z(SUM[14]) );
  XOR2_X1 U115 ( .A(A[6]), .B(n92), .Z(SUM[6]) );
  XOR2_X1 U116 ( .A(A[7]), .B(n93), .Z(SUM[7]) );
  XOR2_X1 U117 ( .A(A[8]), .B(n94), .Z(SUM[8]) );
  XOR2_X1 U118 ( .A(A[9]), .B(n95), .Z(SUM[9]) );
  XOR2_X1 U119 ( .A(A[10]), .B(n78), .Z(SUM[10]) );
  XOR2_X1 U120 ( .A(A[1]), .B(carry[1]), .Z(SUM[1]) );
  XOR2_X1 U121 ( .A(A[2]), .B(n100), .Z(SUM[2]) );
  XOR2_X1 U122 ( .A(A[3]), .B(n89), .Z(SUM[3]) );
  XOR2_X1 U123 ( .A(A[4]), .B(n90), .Z(SUM[4]) );
  XOR2_X1 U124 ( .A(A[5]), .B(n91), .Z(SUM[5]) );
endmodule


module multiplierTreeV2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n11, n23, n24, n25, n26, n27, n28, n29, n31,
         n32, n33, n34, n35, n36, n42, n43, n44, n45, n46, n47, n48, n49;
  wire   [2:1] carry;

  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .S(SUM[0]) );
  FA_X1 U1_1 ( .A(A[1]), .B(1'b0), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(A[5]), .B(n7), .Z(SUM[5]) );
  XOR2_X1 U2 ( .A(A[6]), .B(n8), .Z(SUM[6]) );
  XOR2_X1 U3 ( .A(A[7]), .B(n9), .Z(SUM[7]) );
  XOR2_X1 U4 ( .A(A[8]), .B(n10), .Z(SUM[8]) );
  AND2_X1 U5 ( .A1(A[2]), .A2(carry[2]), .ZN(n5) );
  AND2_X1 U6 ( .A1(A[3]), .A2(n5), .ZN(n6) );
  AND2_X1 U7 ( .A1(A[4]), .A2(n6), .ZN(n7) );
  AND2_X1 U8 ( .A1(A[5]), .A2(n7), .ZN(n8) );
  AND2_X1 U9 ( .A1(A[6]), .A2(n8), .ZN(n9) );
  AND2_X1 U10 ( .A1(A[7]), .A2(n9), .ZN(n10) );
  AND2_X1 U11 ( .A1(A[8]), .A2(n10), .ZN(n11) );
  XOR2_X1 U12 ( .A(A[2]), .B(carry[2]), .Z(SUM[2]) );
  XOR2_X1 U13 ( .A(A[3]), .B(n5), .Z(SUM[3]) );
  XOR2_X1 U14 ( .A(A[4]), .B(n6), .Z(SUM[4]) );
  XOR2_X1 U15 ( .A(A[9]), .B(n11), .Z(SUM[9]) );
  XOR2_X1 U16 ( .A(A[11]), .B(n24), .Z(SUM[11]) );
  XOR2_X1 U17 ( .A(A[12]), .B(n25), .Z(SUM[12]) );
  XOR2_X1 U18 ( .A(A[10]), .B(n23), .Z(SUM[10]) );
  XOR2_X1 U19 ( .A(A[13]), .B(n26), .Z(SUM[13]) );
  XOR2_X1 U20 ( .A(A[14]), .B(n27), .Z(SUM[14]) );
  XOR2_X1 U21 ( .A(A[15]), .B(n28), .Z(SUM[15]) );
  XOR2_X1 U22 ( .A(A[16]), .B(n29), .Z(SUM[16]) );
  AND2_X1 U23 ( .A1(A[9]), .A2(n11), .ZN(n23) );
  AND2_X1 U24 ( .A1(A[10]), .A2(n23), .ZN(n24) );
  AND2_X1 U25 ( .A1(A[11]), .A2(n24), .ZN(n25) );
  AND2_X1 U26 ( .A1(A[12]), .A2(n25), .ZN(n26) );
  AND2_X1 U27 ( .A1(A[13]), .A2(n26), .ZN(n27) );
  AND2_X1 U28 ( .A1(A[14]), .A2(n27), .ZN(n28) );
  AND2_X1 U29 ( .A1(A[15]), .A2(n28), .ZN(n29) );
  XOR2_X1 U30 ( .A(A[17]), .B(n31), .Z(SUM[17]) );
  AND2_X1 U31 ( .A1(A[16]), .A2(n29), .ZN(n31) );
  AND2_X1 U32 ( .A1(A[17]), .A2(n31), .ZN(n32) );
  AND2_X1 U33 ( .A1(A[18]), .A2(n32), .ZN(n33) );
  AND2_X1 U34 ( .A1(A[19]), .A2(n33), .ZN(n34) );
  AND2_X1 U35 ( .A1(A[20]), .A2(n34), .ZN(n35) );
  AND2_X1 U36 ( .A1(A[21]), .A2(n35), .ZN(n36) );
  XOR2_X1 U37 ( .A(A[18]), .B(n32), .Z(SUM[18]) );
  XOR2_X1 U38 ( .A(A[19]), .B(n33), .Z(SUM[19]) );
  XOR2_X1 U39 ( .A(A[20]), .B(n34), .Z(SUM[20]) );
  XOR2_X1 U40 ( .A(A[21]), .B(n35), .Z(SUM[21]) );
  XOR2_X1 U41 ( .A(A[22]), .B(n36), .Z(SUM[22]) );
  AND2_X1 U42 ( .A1(A[22]), .A2(n36), .ZN(n42) );
  AND2_X1 U43 ( .A1(A[23]), .A2(n42), .ZN(n43) );
  AND2_X1 U44 ( .A1(A[24]), .A2(n43), .ZN(n44) );
  AND2_X1 U45 ( .A1(A[25]), .A2(n44), .ZN(n45) );
  AND2_X1 U46 ( .A1(A[26]), .A2(n45), .ZN(n46) );
  AND2_X1 U47 ( .A1(A[27]), .A2(n46), .ZN(n47) );
  AND2_X1 U48 ( .A1(A[28]), .A2(n47), .ZN(n48) );
  AND2_X1 U49 ( .A1(A[29]), .A2(n48), .ZN(n49) );
  XOR2_X1 U50 ( .A(A[24]), .B(n43), .Z(SUM[24]) );
  XOR2_X1 U51 ( .A(A[25]), .B(n44), .Z(SUM[25]) );
  XOR2_X1 U52 ( .A(A[26]), .B(n45), .Z(SUM[26]) );
  XOR2_X1 U53 ( .A(A[27]), .B(n46), .Z(SUM[27]) );
  XOR2_X1 U54 ( .A(A[28]), .B(n47), .Z(SUM[28]) );
  XOR2_X1 U55 ( .A(A[29]), .B(n48), .Z(SUM[29]) );
  XOR2_X1 U56 ( .A(A[30]), .B(n49), .Z(SUM[30]) );
  XOR2_X1 U57 ( .A(A[23]), .B(n42), .Z(SUM[23]) );
  AND2_X1 U58 ( .A1(A[30]), .A2(n49), .ZN(SUM[31]) );
endmodule


module multiplierTreeV2_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n23, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50;

  AND2_X1 U1 ( .A1(A[26]), .A2(n37), .ZN(n1) );
  AND2_X1 U2 ( .A1(A[9]), .A2(n26), .ZN(n2) );
  AND2_X1 U3 ( .A1(A[20]), .A2(n31), .ZN(n3) );
  AND2_X1 U4 ( .A1(A[11]), .A2(n33), .ZN(n39) );
  AND2_X1 U5 ( .A1(A[13]), .A2(n34), .ZN(n40) );
  AND2_X1 U6 ( .A1(A[16]), .A2(n29), .ZN(n41) );
  AND2_X1 U7 ( .A1(A[18]), .A2(n30), .ZN(n42) );
  AND2_X1 U8 ( .A1(A[24]), .A2(n36), .ZN(n44) );
  AND2_X1 U9 ( .A1(A[5]), .A2(n28), .ZN(n47) );
  XOR2_X1 U10 ( .A(A[26]), .B(n37), .Z(SUM[26]) );
  XOR2_X1 U11 ( .A(A[24]), .B(n36), .Z(SUM[24]) );
  XOR2_X1 U12 ( .A(A[14]), .B(n40), .Z(SUM[14]) );
  XOR2_X1 U13 ( .A(A[19]), .B(n42), .Z(SUM[19]) );
  XOR2_X1 U14 ( .A(A[4]), .B(n48), .Z(SUM[4]) );
  XOR2_X1 U15 ( .A(A[29]), .B(n45), .Z(SUM[29]) );
  XOR2_X1 U16 ( .A(A[22]), .B(n32), .Z(SUM[22]) );
  XOR2_X1 U17 ( .A(A[27]), .B(n1), .Z(SUM[27]) );
  XOR2_X1 U18 ( .A(A[25]), .B(n44), .Z(SUM[25]) );
  XOR2_X1 U19 ( .A(A[9]), .B(n26), .Z(SUM[9]) );
  XOR2_X1 U20 ( .A(A[7]), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U21 ( .A(A[21]), .B(n3), .Z(SUM[21]) );
  XOR2_X1 U22 ( .A(A[30]), .B(n46), .Z(SUM[30]) );
  XOR2_X1 U23 ( .A(A[12]), .B(n39), .Z(SUM[12]) );
  XOR2_X1 U24 ( .A(A[10]), .B(n2), .Z(SUM[10]) );
  XOR2_X1 U25 ( .A(A[20]), .B(n31), .Z(SUM[20]) );
  XOR2_X1 U26 ( .A(A[18]), .B(n30), .Z(SUM[18]) );
  XOR2_X1 U27 ( .A(A[23]), .B(n23), .Z(SUM[23]) );
  XOR2_X1 U28 ( .A(A[28]), .B(n38), .Z(SUM[28]) );
  AND2_X1 U29 ( .A1(A[22]), .A2(n32), .ZN(n23) );
  AND2_X1 U30 ( .A1(A[1]), .A2(n50), .ZN(n24) );
  XOR2_X1 U31 ( .A(A[15]), .B(n35), .Z(SUM[15]) );
  AND2_X1 U32 ( .A1(A[8]), .A2(n43), .ZN(n26) );
  AND2_X1 U33 ( .A1(A[6]), .A2(n47), .ZN(n27) );
  AND2_X1 U34 ( .A1(A[4]), .A2(n48), .ZN(n28) );
  AND2_X1 U35 ( .A1(A[15]), .A2(n35), .ZN(n29) );
  AND2_X1 U36 ( .A1(A[17]), .A2(n41), .ZN(n30) );
  AND2_X1 U37 ( .A1(A[19]), .A2(n42), .ZN(n31) );
  AND2_X1 U38 ( .A1(A[21]), .A2(n3), .ZN(n32) );
  AND2_X1 U39 ( .A1(A[10]), .A2(n2), .ZN(n33) );
  AND2_X1 U40 ( .A1(A[12]), .A2(n39), .ZN(n34) );
  AND2_X1 U41 ( .A1(A[14]), .A2(n40), .ZN(n35) );
  AND2_X1 U42 ( .A1(A[23]), .A2(n23), .ZN(n36) );
  AND2_X1 U43 ( .A1(A[25]), .A2(n44), .ZN(n37) );
  AND2_X1 U44 ( .A1(A[27]), .A2(n1), .ZN(n38) );
  AND2_X1 U45 ( .A1(A[7]), .A2(n27), .ZN(n43) );
  AND2_X1 U46 ( .A1(A[28]), .A2(n38), .ZN(n45) );
  AND2_X1 U47 ( .A1(A[29]), .A2(n45), .ZN(n46) );
  AND2_X1 U48 ( .A1(A[3]), .A2(n49), .ZN(n48) );
  AND2_X1 U49 ( .A1(A[2]), .A2(n24), .ZN(n49) );
  AND2_X1 U50 ( .A1(B[0]), .A2(A[0]), .ZN(n50) );
  XOR2_X1 U51 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  XOR2_X1 U52 ( .A(A[17]), .B(n41), .Z(SUM[17]) );
  XOR2_X1 U53 ( .A(A[8]), .B(n43), .Z(SUM[8]) );
  XOR2_X1 U54 ( .A(A[16]), .B(n29), .Z(SUM[16]) );
  XOR2_X1 U55 ( .A(A[13]), .B(n34), .Z(SUM[13]) );
  XOR2_X1 U56 ( .A(A[3]), .B(n49), .Z(SUM[3]) );
  XOR2_X1 U57 ( .A(A[5]), .B(n28), .Z(SUM[5]) );
  XOR2_X1 U58 ( .A(A[2]), .B(n24), .Z(SUM[2]) );
  XOR2_X1 U59 ( .A(A[1]), .B(n50), .Z(SUM[1]) );
  AND2_X1 U60 ( .A1(A[30]), .A2(n46), .ZN(SUM[31]) );
  XOR2_X1 U61 ( .A(A[6]), .B(n47), .Z(SUM[6]) );
  XOR2_X1 U62 ( .A(A[11]), .B(n33), .Z(SUM[11]) );
endmodule


module multiplierTreeV2 ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, finalSign, tempResultA_30__31_,
         tempResultA_30__30_, tempResultA_30__29_, tempResultA_30__28_,
         tempResultA_30__27_, tempResultA_30__26_, tempResultA_30__25_,
         tempResultA_30__24_, tempResultA_30__23_, tempResultA_30__22_,
         tempResultA_30__21_, tempResultA_30__20_, tempResultA_30__19_,
         tempResultA_30__18_, tempResultA_30__17_, tempResultA_30__16_,
         tempResultA_30__15_, tempResultA_30__14_, tempResultA_30__13_,
         tempResultA_30__12_, tempResultA_30__11_, tempResultA_30__10_,
         tempResultA_30__9_, tempResultA_30__8_, tempResultA_30__7_,
         tempResultA_30__6_, tempResultA_30__5_, tempResultA_30__4_,
         tempResultA_30__3_, tempResultA_30__2_, tempResultA_30__1_,
         tempResultA_30__0_, tempResultA_29__31_, tempResultA_29__30_,
         tempResultA_29__29_, tempResultA_29__28_, tempResultA_29__27_,
         tempResultA_29__26_, tempResultA_29__25_, tempResultA_29__24_,
         tempResultA_29__23_, tempResultA_29__22_, tempResultA_29__21_,
         tempResultA_29__20_, tempResultA_29__19_, tempResultA_29__18_,
         tempResultA_29__17_, tempResultA_29__16_, tempResultA_29__15_,
         tempResultA_29__14_, tempResultA_29__13_, tempResultA_29__12_,
         tempResultA_29__11_, tempResultA_29__10_, tempResultA_29__9_,
         tempResultA_29__8_, tempResultA_29__7_, tempResultA_29__6_,
         tempResultA_29__5_, tempResultA_29__4_, tempResultA_29__3_,
         tempResultA_29__2_, tempResultA_29__1_, tempResultA_29__0_,
         tempResultA_28__31_, tempResultA_28__30_, tempResultA_28__29_,
         tempResultA_28__28_, tempResultA_28__27_, tempResultA_28__26_,
         tempResultA_28__25_, tempResultA_28__24_, tempResultA_28__23_,
         tempResultA_28__22_, tempResultA_28__21_, tempResultA_28__20_,
         tempResultA_28__19_, tempResultA_28__18_, tempResultA_28__17_,
         tempResultA_28__16_, tempResultA_28__15_, tempResultA_28__14_,
         tempResultA_28__13_, tempResultA_28__12_, tempResultA_28__11_,
         tempResultA_28__10_, tempResultA_28__9_, tempResultA_28__8_,
         tempResultA_28__7_, tempResultA_28__6_, tempResultA_28__5_,
         tempResultA_28__4_, tempResultA_28__3_, tempResultA_28__2_,
         tempResultA_28__1_, tempResultA_28__0_, tempResultA_27__31_,
         tempResultA_27__30_, tempResultA_27__29_, tempResultA_27__28_,
         tempResultA_27__27_, tempResultA_27__26_, tempResultA_27__25_,
         tempResultA_27__24_, tempResultA_27__23_, tempResultA_27__22_,
         tempResultA_27__21_, tempResultA_27__20_, tempResultA_27__19_,
         tempResultA_27__18_, tempResultA_27__17_, tempResultA_27__16_,
         tempResultA_27__15_, tempResultA_27__14_, tempResultA_27__13_,
         tempResultA_27__12_, tempResultA_27__11_, tempResultA_27__10_,
         tempResultA_27__9_, tempResultA_27__8_, tempResultA_27__7_,
         tempResultA_27__6_, tempResultA_27__5_, tempResultA_27__4_,
         tempResultA_27__3_, tempResultA_27__2_, tempResultA_27__1_,
         tempResultA_27__0_, tempResultA_26__31_, tempResultA_26__30_,
         tempResultA_26__29_, tempResultA_26__28_, tempResultA_26__27_,
         tempResultA_26__26_, tempResultA_26__25_, tempResultA_26__24_,
         tempResultA_26__23_, tempResultA_26__22_, tempResultA_26__21_,
         tempResultA_26__20_, tempResultA_26__19_, tempResultA_26__18_,
         tempResultA_26__17_, tempResultA_26__16_, tempResultA_26__15_,
         tempResultA_26__14_, tempResultA_26__13_, tempResultA_26__12_,
         tempResultA_26__11_, tempResultA_26__10_, tempResultA_26__9_,
         tempResultA_26__8_, tempResultA_26__7_, tempResultA_26__6_,
         tempResultA_26__5_, tempResultA_26__4_, tempResultA_26__3_,
         tempResultA_26__2_, tempResultA_26__1_, tempResultA_26__0_,
         tempResultA_25__31_, tempResultA_25__30_, tempResultA_25__29_,
         tempResultA_25__28_, tempResultA_25__27_, tempResultA_25__26_,
         tempResultA_25__25_, tempResultA_25__24_, tempResultA_25__23_,
         tempResultA_25__22_, tempResultA_25__21_, tempResultA_25__20_,
         tempResultA_25__19_, tempResultA_25__18_, tempResultA_25__17_,
         tempResultA_25__16_, tempResultA_25__15_, tempResultA_25__14_,
         tempResultA_25__13_, tempResultA_25__12_, tempResultA_25__11_,
         tempResultA_25__10_, tempResultA_25__9_, tempResultA_25__8_,
         tempResultA_25__7_, tempResultA_25__6_, tempResultA_25__5_,
         tempResultA_25__4_, tempResultA_25__3_, tempResultA_25__2_,
         tempResultA_25__1_, tempResultA_25__0_, tempResultA_24__31_,
         tempResultA_24__30_, tempResultA_24__29_, tempResultA_24__28_,
         tempResultA_24__27_, tempResultA_24__26_, tempResultA_24__25_,
         tempResultA_24__24_, tempResultA_24__23_, tempResultA_24__22_,
         tempResultA_24__21_, tempResultA_24__20_, tempResultA_24__19_,
         tempResultA_24__18_, tempResultA_24__17_, tempResultA_24__16_,
         tempResultA_24__15_, tempResultA_24__14_, tempResultA_24__13_,
         tempResultA_24__12_, tempResultA_24__11_, tempResultA_24__10_,
         tempResultA_24__9_, tempResultA_24__8_, tempResultA_24__7_,
         tempResultA_24__6_, tempResultA_24__5_, tempResultA_24__4_,
         tempResultA_24__3_, tempResultA_24__2_, tempResultA_24__1_,
         tempResultA_24__0_, tempResultA_23__31_, tempResultA_23__30_,
         tempResultA_23__29_, tempResultA_23__28_, tempResultA_23__27_,
         tempResultA_23__26_, tempResultA_23__25_, tempResultA_23__24_,
         tempResultA_23__23_, tempResultA_23__22_, tempResultA_23__21_,
         tempResultA_23__20_, tempResultA_23__19_, tempResultA_23__18_,
         tempResultA_23__17_, tempResultA_23__16_, tempResultA_23__15_,
         tempResultA_23__14_, tempResultA_23__13_, tempResultA_23__12_,
         tempResultA_23__11_, tempResultA_23__10_, tempResultA_23__9_,
         tempResultA_23__8_, tempResultA_23__7_, tempResultA_23__6_,
         tempResultA_23__5_, tempResultA_23__4_, tempResultA_23__3_,
         tempResultA_23__2_, tempResultA_23__1_, tempResultA_23__0_,
         tempResultA_22__31_, tempResultA_22__30_, tempResultA_22__29_,
         tempResultA_22__28_, tempResultA_22__27_, tempResultA_22__26_,
         tempResultA_22__25_, tempResultA_22__24_, tempResultA_22__23_,
         tempResultA_22__22_, tempResultA_22__21_, tempResultA_22__20_,
         tempResultA_22__19_, tempResultA_22__18_, tempResultA_22__17_,
         tempResultA_22__16_, tempResultA_22__15_, tempResultA_22__14_,
         tempResultA_22__13_, tempResultA_22__12_, tempResultA_22__11_,
         tempResultA_22__10_, tempResultA_22__9_, tempResultA_22__8_,
         tempResultA_22__7_, tempResultA_22__6_, tempResultA_22__5_,
         tempResultA_22__4_, tempResultA_22__3_, tempResultA_22__2_,
         tempResultA_22__1_, tempResultA_22__0_, tempResultA_21__31_,
         tempResultA_21__30_, tempResultA_21__29_, tempResultA_21__28_,
         tempResultA_21__27_, tempResultA_21__26_, tempResultA_21__25_,
         tempResultA_21__24_, tempResultA_21__23_, tempResultA_21__22_,
         tempResultA_21__21_, tempResultA_21__20_, tempResultA_21__19_,
         tempResultA_21__18_, tempResultA_21__17_, tempResultA_21__16_,
         tempResultA_21__15_, tempResultA_21__14_, tempResultA_21__13_,
         tempResultA_21__12_, tempResultA_21__11_, tempResultA_21__10_,
         tempResultA_21__9_, tempResultA_21__8_, tempResultA_21__7_,
         tempResultA_21__6_, tempResultA_21__5_, tempResultA_21__4_,
         tempResultA_21__3_, tempResultA_21__2_, tempResultA_21__1_,
         tempResultA_21__0_, tempResultA_20__31_, tempResultA_20__30_,
         tempResultA_20__29_, tempResultA_20__28_, tempResultA_20__27_,
         tempResultA_20__26_, tempResultA_20__25_, tempResultA_20__24_,
         tempResultA_20__23_, tempResultA_20__22_, tempResultA_20__21_,
         tempResultA_20__20_, tempResultA_20__19_, tempResultA_20__18_,
         tempResultA_20__17_, tempResultA_20__16_, tempResultA_20__15_,
         tempResultA_20__14_, tempResultA_20__13_, tempResultA_20__12_,
         tempResultA_20__11_, tempResultA_20__10_, tempResultA_20__9_,
         tempResultA_20__8_, tempResultA_20__7_, tempResultA_20__6_,
         tempResultA_20__5_, tempResultA_20__4_, tempResultA_20__3_,
         tempResultA_20__2_, tempResultA_20__1_, tempResultA_20__0_,
         tempResultA_19__31_, tempResultA_19__30_, tempResultA_19__29_,
         tempResultA_19__28_, tempResultA_19__27_, tempResultA_19__26_,
         tempResultA_19__25_, tempResultA_19__24_, tempResultA_19__23_,
         tempResultA_19__22_, tempResultA_19__21_, tempResultA_19__20_,
         tempResultA_19__19_, tempResultA_19__18_, tempResultA_19__17_,
         tempResultA_19__16_, tempResultA_19__15_, tempResultA_19__14_,
         tempResultA_19__13_, tempResultA_19__12_, tempResultA_19__11_,
         tempResultA_19__10_, tempResultA_19__9_, tempResultA_19__8_,
         tempResultA_19__7_, tempResultA_19__6_, tempResultA_19__5_,
         tempResultA_19__4_, tempResultA_19__3_, tempResultA_19__2_,
         tempResultA_19__1_, tempResultA_19__0_, tempResultA_18__31_,
         tempResultA_18__30_, tempResultA_18__29_, tempResultA_18__28_,
         tempResultA_18__27_, tempResultA_18__26_, tempResultA_18__25_,
         tempResultA_18__24_, tempResultA_18__23_, tempResultA_18__22_,
         tempResultA_18__21_, tempResultA_18__20_, tempResultA_18__19_,
         tempResultA_18__18_, tempResultA_18__17_, tempResultA_18__16_,
         tempResultA_18__15_, tempResultA_18__14_, tempResultA_18__13_,
         tempResultA_18__12_, tempResultA_18__11_, tempResultA_18__10_,
         tempResultA_18__9_, tempResultA_18__8_, tempResultA_18__7_,
         tempResultA_18__6_, tempResultA_18__5_, tempResultA_18__4_,
         tempResultA_18__3_, tempResultA_18__2_, tempResultA_18__1_,
         tempResultA_18__0_, tempResultA_17__31_, tempResultA_17__30_,
         tempResultA_17__29_, tempResultA_17__28_, tempResultA_17__27_,
         tempResultA_17__26_, tempResultA_17__25_, tempResultA_17__24_,
         tempResultA_17__23_, tempResultA_17__22_, tempResultA_17__21_,
         tempResultA_17__20_, tempResultA_17__19_, tempResultA_17__18_,
         tempResultA_17__17_, tempResultA_17__16_, tempResultA_17__15_,
         tempResultA_17__14_, tempResultA_17__13_, tempResultA_17__12_,
         tempResultA_17__11_, tempResultA_17__10_, tempResultA_17__9_,
         tempResultA_17__8_, tempResultA_17__7_, tempResultA_17__6_,
         tempResultA_17__5_, tempResultA_17__4_, tempResultA_17__3_,
         tempResultA_17__2_, tempResultA_17__1_, tempResultA_17__0_,
         tempResultA_16__31_, tempResultA_16__30_, tempResultA_16__29_,
         tempResultA_16__28_, tempResultA_16__27_, tempResultA_16__26_,
         tempResultA_16__25_, tempResultA_16__24_, tempResultA_16__23_,
         tempResultA_16__22_, tempResultA_16__21_, tempResultA_16__20_,
         tempResultA_16__19_, tempResultA_16__18_, tempResultA_16__17_,
         tempResultA_16__16_, tempResultA_16__15_, tempResultA_16__14_,
         tempResultA_16__13_, tempResultA_16__12_, tempResultA_16__11_,
         tempResultA_16__10_, tempResultA_16__9_, tempResultA_16__8_,
         tempResultA_16__7_, tempResultA_16__6_, tempResultA_16__5_,
         tempResultA_16__4_, tempResultA_16__3_, tempResultA_16__2_,
         tempResultA_16__1_, tempResultA_16__0_, tempResultA_15__31_,
         tempResultA_15__30_, tempResultA_15__29_, tempResultA_15__28_,
         tempResultA_15__27_, tempResultA_15__26_, tempResultA_15__25_,
         tempResultA_15__24_, tempResultA_15__23_, tempResultA_15__22_,
         tempResultA_15__21_, tempResultA_15__20_, tempResultA_15__19_,
         tempResultA_15__18_, tempResultA_15__17_, tempResultA_15__16_,
         tempResultA_15__15_, tempResultA_15__14_, tempResultA_15__13_,
         tempResultA_15__12_, tempResultA_15__11_, tempResultA_15__10_,
         tempResultA_15__9_, tempResultA_15__8_, tempResultA_15__7_,
         tempResultA_15__6_, tempResultA_15__5_, tempResultA_15__4_,
         tempResultA_15__3_, tempResultA_15__2_, tempResultA_15__1_,
         tempResultA_15__0_, tempResultA_14__31_, tempResultA_14__30_,
         tempResultA_14__29_, tempResultA_14__28_, tempResultA_14__27_,
         tempResultA_14__26_, tempResultA_14__25_, tempResultA_14__24_,
         tempResultA_14__23_, tempResultA_14__22_, tempResultA_14__21_,
         tempResultA_14__20_, tempResultA_14__19_, tempResultA_14__18_,
         tempResultA_14__17_, tempResultA_14__16_, tempResultA_14__15_,
         tempResultA_14__14_, tempResultA_14__13_, tempResultA_14__12_,
         tempResultA_14__11_, tempResultA_14__10_, tempResultA_14__9_,
         tempResultA_14__8_, tempResultA_14__7_, tempResultA_14__6_,
         tempResultA_14__5_, tempResultA_14__4_, tempResultA_14__3_,
         tempResultA_14__2_, tempResultA_14__1_, tempResultA_14__0_,
         tempResultA_13__31_, tempResultA_13__30_, tempResultA_13__29_,
         tempResultA_13__28_, tempResultA_13__27_, tempResultA_13__26_,
         tempResultA_13__25_, tempResultA_13__24_, tempResultA_13__23_,
         tempResultA_13__22_, tempResultA_13__21_, tempResultA_13__20_,
         tempResultA_13__19_, tempResultA_13__18_, tempResultA_13__17_,
         tempResultA_13__16_, tempResultA_13__15_, tempResultA_13__14_,
         tempResultA_13__13_, tempResultA_13__12_, tempResultA_13__11_,
         tempResultA_13__10_, tempResultA_13__9_, tempResultA_13__8_,
         tempResultA_13__7_, tempResultA_13__6_, tempResultA_13__5_,
         tempResultA_13__4_, tempResultA_13__3_, tempResultA_13__2_,
         tempResultA_13__1_, tempResultA_13__0_, tempResultA_12__31_,
         tempResultA_12__30_, tempResultA_12__29_, tempResultA_12__28_,
         tempResultA_12__27_, tempResultA_12__26_, tempResultA_12__25_,
         tempResultA_12__24_, tempResultA_12__23_, tempResultA_12__22_,
         tempResultA_12__21_, tempResultA_12__20_, tempResultA_12__19_,
         tempResultA_12__18_, tempResultA_12__17_, tempResultA_12__16_,
         tempResultA_12__15_, tempResultA_12__14_, tempResultA_12__13_,
         tempResultA_12__12_, tempResultA_12__11_, tempResultA_12__10_,
         tempResultA_12__9_, tempResultA_12__8_, tempResultA_12__7_,
         tempResultA_12__6_, tempResultA_12__5_, tempResultA_12__4_,
         tempResultA_12__3_, tempResultA_12__2_, tempResultA_12__1_,
         tempResultA_12__0_, tempResultA_11__31_, tempResultA_11__30_,
         tempResultA_11__29_, tempResultA_11__28_, tempResultA_11__27_,
         tempResultA_11__26_, tempResultA_11__25_, tempResultA_11__24_,
         tempResultA_11__23_, tempResultA_11__22_, tempResultA_11__21_,
         tempResultA_11__20_, tempResultA_11__19_, tempResultA_11__18_,
         tempResultA_11__17_, tempResultA_11__16_, tempResultA_11__15_,
         tempResultA_11__14_, tempResultA_11__13_, tempResultA_11__12_,
         tempResultA_11__11_, tempResultA_11__10_, tempResultA_11__9_,
         tempResultA_11__8_, tempResultA_11__7_, tempResultA_11__6_,
         tempResultA_11__5_, tempResultA_11__4_, tempResultA_11__3_,
         tempResultA_11__2_, tempResultA_11__1_, tempResultA_11__0_,
         tempResultA_10__31_, tempResultA_10__30_, tempResultA_10__29_,
         tempResultA_10__28_, tempResultA_10__27_, tempResultA_10__26_,
         tempResultA_10__25_, tempResultA_10__24_, tempResultA_10__23_,
         tempResultA_10__22_, tempResultA_10__21_, tempResultA_10__20_,
         tempResultA_10__19_, tempResultA_10__18_, tempResultA_10__17_,
         tempResultA_10__16_, tempResultA_10__15_, tempResultA_10__14_,
         tempResultA_10__13_, tempResultA_10__12_, tempResultA_10__11_,
         tempResultA_10__10_, tempResultA_10__9_, tempResultA_10__8_,
         tempResultA_10__7_, tempResultA_10__6_, tempResultA_10__5_,
         tempResultA_10__4_, tempResultA_10__3_, tempResultA_10__2_,
         tempResultA_10__1_, tempResultA_10__0_, tempResultA_9__31_,
         tempResultA_9__30_, tempResultA_9__29_, tempResultA_9__28_,
         tempResultA_9__27_, tempResultA_9__26_, tempResultA_9__25_,
         tempResultA_9__24_, tempResultA_9__23_, tempResultA_9__22_,
         tempResultA_9__21_, tempResultA_9__20_, tempResultA_9__19_,
         tempResultA_9__18_, tempResultA_9__17_, tempResultA_9__16_,
         tempResultA_9__15_, tempResultA_9__14_, tempResultA_9__13_,
         tempResultA_9__12_, tempResultA_9__11_, tempResultA_9__10_,
         tempResultA_9__9_, tempResultA_9__8_, tempResultA_9__7_,
         tempResultA_9__6_, tempResultA_9__5_, tempResultA_9__4_,
         tempResultA_9__3_, tempResultA_9__2_, tempResultA_9__1_,
         tempResultA_9__0_, tempResultA_8__31_, tempResultA_8__30_,
         tempResultA_8__29_, tempResultA_8__28_, tempResultA_8__27_,
         tempResultA_8__26_, tempResultA_8__25_, tempResultA_8__24_,
         tempResultA_8__23_, tempResultA_8__22_, tempResultA_8__21_,
         tempResultA_8__20_, tempResultA_8__19_, tempResultA_8__18_,
         tempResultA_8__17_, tempResultA_8__16_, tempResultA_8__15_,
         tempResultA_8__14_, tempResultA_8__13_, tempResultA_8__12_,
         tempResultA_8__11_, tempResultA_8__10_, tempResultA_8__9_,
         tempResultA_8__8_, tempResultA_8__7_, tempResultA_8__6_,
         tempResultA_8__5_, tempResultA_8__4_, tempResultA_8__3_,
         tempResultA_8__2_, tempResultA_8__1_, tempResultA_8__0_,
         tempResultA_7__31_, tempResultA_7__30_, tempResultA_7__29_,
         tempResultA_7__28_, tempResultA_7__27_, tempResultA_7__26_,
         tempResultA_7__25_, tempResultA_7__24_, tempResultA_7__23_,
         tempResultA_7__22_, tempResultA_7__21_, tempResultA_7__20_,
         tempResultA_7__19_, tempResultA_7__18_, tempResultA_7__17_,
         tempResultA_7__16_, tempResultA_7__15_, tempResultA_7__14_,
         tempResultA_7__13_, tempResultA_7__12_, tempResultA_7__11_,
         tempResultA_7__10_, tempResultA_7__9_, tempResultA_7__8_,
         tempResultA_7__7_, tempResultA_7__6_, tempResultA_7__5_,
         tempResultA_7__4_, tempResultA_7__3_, tempResultA_7__2_,
         tempResultA_7__1_, tempResultA_7__0_, tempResultA_6__31_,
         tempResultA_6__30_, tempResultA_6__29_, tempResultA_6__28_,
         tempResultA_6__27_, tempResultA_6__26_, tempResultA_6__25_,
         tempResultA_6__24_, tempResultA_6__23_, tempResultA_6__22_,
         tempResultA_6__21_, tempResultA_6__20_, tempResultA_6__19_,
         tempResultA_6__18_, tempResultA_6__17_, tempResultA_6__16_,
         tempResultA_6__15_, tempResultA_6__14_, tempResultA_6__13_,
         tempResultA_6__12_, tempResultA_6__11_, tempResultA_6__10_,
         tempResultA_6__9_, tempResultA_6__8_, tempResultA_6__7_,
         tempResultA_6__6_, tempResultA_6__5_, tempResultA_6__4_,
         tempResultA_6__3_, tempResultA_6__2_, tempResultA_6__1_,
         tempResultA_6__0_, tempResultA_5__31_, tempResultA_5__30_,
         tempResultA_5__29_, tempResultA_5__28_, tempResultA_5__27_,
         tempResultA_5__26_, tempResultA_5__25_, tempResultA_5__24_,
         tempResultA_5__23_, tempResultA_5__22_, tempResultA_5__21_,
         tempResultA_5__20_, tempResultA_5__19_, tempResultA_5__18_,
         tempResultA_5__17_, tempResultA_5__16_, tempResultA_5__15_,
         tempResultA_5__14_, tempResultA_5__13_, tempResultA_5__12_,
         tempResultA_5__11_, tempResultA_5__10_, tempResultA_5__9_,
         tempResultA_5__8_, tempResultA_5__7_, tempResultA_5__6_,
         tempResultA_5__5_, tempResultA_5__4_, tempResultA_5__3_,
         tempResultA_5__2_, tempResultA_5__1_, tempResultA_5__0_,
         tempResultA_4__31_, tempResultA_4__30_, tempResultA_4__29_,
         tempResultA_4__28_, tempResultA_4__27_, tempResultA_4__26_,
         tempResultA_4__25_, tempResultA_4__24_, tempResultA_4__23_,
         tempResultA_4__22_, tempResultA_4__21_, tempResultA_4__20_,
         tempResultA_4__19_, tempResultA_4__18_, tempResultA_4__17_,
         tempResultA_4__16_, tempResultA_4__15_, tempResultA_4__14_,
         tempResultA_4__13_, tempResultA_4__12_, tempResultA_4__11_,
         tempResultA_4__10_, tempResultA_4__9_, tempResultA_4__8_,
         tempResultA_4__7_, tempResultA_4__6_, tempResultA_4__5_,
         tempResultA_4__4_, tempResultA_4__3_, tempResultA_4__2_,
         tempResultA_4__1_, tempResultA_4__0_, tempResultA_3__31_,
         tempResultA_3__30_, tempResultA_3__29_, tempResultA_3__28_,
         tempResultA_3__27_, tempResultA_3__26_, tempResultA_3__25_,
         tempResultA_3__24_, tempResultA_3__23_, tempResultA_3__22_,
         tempResultA_3__21_, tempResultA_3__20_, tempResultA_3__19_,
         tempResultA_3__18_, tempResultA_3__17_, tempResultA_3__16_,
         tempResultA_3__15_, tempResultA_3__14_, tempResultA_3__13_,
         tempResultA_3__12_, tempResultA_3__11_, tempResultA_3__10_,
         tempResultA_3__9_, tempResultA_3__8_, tempResultA_3__7_,
         tempResultA_3__6_, tempResultA_3__5_, tempResultA_3__4_,
         tempResultA_3__3_, tempResultA_3__2_, tempResultA_3__1_,
         tempResultA_3__0_, tempResultA_2__31_, tempResultA_2__30_,
         tempResultA_2__29_, tempResultA_2__28_, tempResultA_2__27_,
         tempResultA_2__26_, tempResultA_2__25_, tempResultA_2__24_,
         tempResultA_2__23_, tempResultA_2__22_, tempResultA_2__21_,
         tempResultA_2__20_, tempResultA_2__19_, tempResultA_2__18_,
         tempResultA_2__17_, tempResultA_2__16_, tempResultA_2__15_,
         tempResultA_2__14_, tempResultA_2__13_, tempResultA_2__12_,
         tempResultA_2__11_, tempResultA_2__10_, tempResultA_2__9_,
         tempResultA_2__8_, tempResultA_2__7_, tempResultA_2__6_,
         tempResultA_2__5_, tempResultA_2__4_, tempResultA_2__3_,
         tempResultA_2__2_, tempResultA_2__1_, tempResultA_2__0_,
         tempResultA_1__31_, tempResultA_1__30_, tempResultA_1__29_,
         tempResultA_1__28_, tempResultA_1__27_, tempResultA_1__26_,
         tempResultA_1__25_, tempResultA_1__24_, tempResultA_1__23_,
         tempResultA_1__22_, tempResultA_1__21_, tempResultA_1__20_,
         tempResultA_1__19_, tempResultA_1__18_, tempResultA_1__17_,
         tempResultA_1__16_, tempResultA_1__15_, tempResultA_1__14_,
         tempResultA_1__13_, tempResultA_1__12_, tempResultA_1__11_,
         tempResultA_1__10_, tempResultA_1__9_, tempResultA_1__8_,
         tempResultA_1__7_, tempResultA_1__6_, tempResultA_1__5_,
         tempResultA_1__4_, tempResultA_1__3_, tempResultA_1__2_,
         tempResultA_1__1_, tempResultA_1__0_, tempResultA_0__30_,
         tempResultA_0__29_, tempResultA_0__28_, tempResultA_0__27_,
         tempResultA_0__26_, tempResultA_0__25_, tempResultA_0__24_,
         tempResultA_0__23_, tempResultA_0__22_, tempResultA_0__21_,
         tempResultA_0__20_, tempResultA_0__19_, tempResultA_0__18_,
         tempResultA_0__17_, tempResultA_0__16_, tempResultA_0__15_,
         tempResultA_0__14_, tempResultA_0__13_, tempResultA_0__12_,
         tempResultA_0__11_, tempResultA_0__10_, tempResultA_0__9_,
         tempResultA_0__8_, tempResultA_0__7_, tempResultA_0__6_,
         tempResultA_0__5_, tempResultA_0__4_, tempResultA_0__3_,
         tempResultA_0__2_, tempResultA_0__1_, tempResultA_0__0_, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104,
         N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115,
         N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, n68, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263;
  wire   [31:0] a_abs;
  wire   [31:0] b_abs;
  wire   [991:0] tempResultB;
  wire   [63:1] tempResult;

  XOR2_X1 U1093 ( .A(tempResult[26]), .B(n193), .Z(N99) );
  XOR2_X1 U1094 ( .A(tempResult[27]), .B(n193), .Z(N98) );
  XOR2_X1 U1095 ( .A(tempResult[28]), .B(n193), .Z(N97) );
  XOR2_X1 U1096 ( .A(tempResult[29]), .B(n193), .Z(N96) );
  XOR2_X1 U1097 ( .A(tempResult[30]), .B(n193), .Z(N95) );
  XOR2_X1 U1098 ( .A(tempResult[31]), .B(n193), .Z(N94) );
  XOR2_X1 U1099 ( .A(tempResult[32]), .B(n193), .Z(N93) );
  XOR2_X1 U1100 ( .A(tempResult[33]), .B(n193), .Z(N92) );
  XOR2_X1 U1102 ( .A(tempResult[35]), .B(n193), .Z(N90) );
  XOR2_X1 U1103 ( .A(n6), .B(a[21]), .Z(N9) );
  XOR2_X1 U1104 ( .A(tempResult[36]), .B(n193), .Z(N89) );
  XOR2_X1 U1105 ( .A(tempResult[37]), .B(n193), .Z(N88) );
  XOR2_X1 U1106 ( .A(tempResult[38]), .B(n193), .Z(N87) );
  XOR2_X1 U1107 ( .A(tempResult[39]), .B(n193), .Z(N86) );
  XOR2_X1 U1108 ( .A(tempResult[40]), .B(n193), .Z(N85) );
  XOR2_X1 U1109 ( .A(tempResult[41]), .B(n193), .Z(N84) );
  XOR2_X1 U1110 ( .A(tempResult[42]), .B(n194), .Z(N83) );
  XOR2_X1 U1111 ( .A(tempResult[43]), .B(n194), .Z(N82) );
  XOR2_X1 U1112 ( .A(tempResult[44]), .B(n194), .Z(N81) );
  XOR2_X1 U1113 ( .A(tempResult[45]), .B(n194), .Z(N80) );
  XOR2_X1 U1114 ( .A(n5), .B(a[22]), .Z(N8) );
  XOR2_X1 U1115 ( .A(tempResult[46]), .B(n194), .Z(N79) );
  XOR2_X1 U1116 ( .A(tempResult[47]), .B(n194), .Z(N78) );
  XOR2_X1 U1117 ( .A(tempResult[48]), .B(n194), .Z(N77) );
  XOR2_X1 U1118 ( .A(tempResult[49]), .B(n194), .Z(N76) );
  XOR2_X1 U1119 ( .A(tempResult[50]), .B(n194), .Z(N75) );
  XOR2_X1 U1120 ( .A(tempResult[51]), .B(n194), .Z(N74) );
  XOR2_X1 U1121 ( .A(tempResult[52]), .B(n194), .Z(N73) );
  XOR2_X1 U1122 ( .A(tempResult[53]), .B(n194), .Z(N72) );
  XOR2_X1 U1123 ( .A(tempResult[54]), .B(n194), .Z(N71) );
  XOR2_X1 U1124 ( .A(tempResult[55]), .B(n194), .Z(N70) );
  XOR2_X1 U1125 ( .A(n4), .B(a[23]), .Z(N7) );
  XOR2_X1 U1126 ( .A(tempResult[56]), .B(n194), .Z(N69) );
  XOR2_X1 U1127 ( .A(tempResult[57]), .B(n194), .Z(N68) );
  XOR2_X1 U1128 ( .A(tempResult[58]), .B(n194), .Z(N67) );
  XOR2_X1 U1129 ( .A(tempResult[59]), .B(n195), .Z(N66) );
  XOR2_X1 U1130 ( .A(tempResult[60]), .B(n195), .Z(N65) );
  XOR2_X1 U1131 ( .A(tempResult[61]), .B(n195), .Z(N64) );
  XOR2_X1 U1132 ( .A(tempResult[62]), .B(n195), .Z(N63) );
  XOR2_X1 U1133 ( .A(tempResult[63]), .B(n195), .Z(N62) );
  XOR2_X1 U1134 ( .A(b[31]), .B(b[0]), .Z(N61) );
  XOR2_X1 U1135 ( .A(n198), .B(b[1]), .Z(N60) );
  XOR2_X1 U1136 ( .A(n5), .B(a[24]), .Z(N6) );
  XOR2_X1 U1137 ( .A(n198), .B(b[2]), .Z(N59) );
  XOR2_X1 U1138 ( .A(b[3]), .B(n197), .Z(N58) );
  XOR2_X1 U1139 ( .A(b[4]), .B(n197), .Z(N57) );
  XOR2_X1 U1140 ( .A(b[5]), .B(n197), .Z(N56) );
  XOR2_X1 U1141 ( .A(b[6]), .B(n197), .Z(N55) );
  XOR2_X1 U1142 ( .A(b[7]), .B(n197), .Z(N54) );
  XOR2_X1 U1143 ( .A(b[8]), .B(n197), .Z(N53) );
  XOR2_X1 U1144 ( .A(b[9]), .B(n197), .Z(N52) );
  XOR2_X1 U1145 ( .A(n198), .B(b[10]), .Z(N51) );
  XOR2_X1 U1146 ( .A(n198), .B(b[11]), .Z(N50) );
  XOR2_X1 U1147 ( .A(n4), .B(a[25]), .Z(N5) );
  XOR2_X1 U1148 ( .A(n198), .B(b[12]), .Z(N49) );
  XOR2_X1 U1149 ( .A(n198), .B(b[13]), .Z(N48) );
  XOR2_X1 U1150 ( .A(n198), .B(b[14]), .Z(N47) );
  XOR2_X1 U1151 ( .A(n198), .B(b[15]), .Z(N46) );
  XOR2_X1 U1152 ( .A(n198), .B(b[16]), .Z(N45) );
  XOR2_X1 U1153 ( .A(n198), .B(b[17]), .Z(N44) );
  XOR2_X1 U1154 ( .A(n198), .B(b[18]), .Z(N43) );
  XOR2_X1 U1155 ( .A(n198), .B(b[19]), .Z(N42) );
  XOR2_X1 U1156 ( .A(n198), .B(b[20]), .Z(N41) );
  XOR2_X1 U1157 ( .A(n198), .B(b[21]), .Z(N40) );
  XOR2_X1 U1158 ( .A(n5), .B(a[26]), .Z(N4) );
  XOR2_X1 U1159 ( .A(n198), .B(b[22]), .Z(N39) );
  XOR2_X1 U1160 ( .A(n198), .B(b[23]), .Z(N38) );
  XOR2_X1 U1161 ( .A(n197), .B(b[24]), .Z(N37) );
  XOR2_X1 U1162 ( .A(n197), .B(b[25]), .Z(N36) );
  XOR2_X1 U1163 ( .A(n197), .B(b[26]), .Z(N35) );
  XOR2_X1 U1164 ( .A(n197), .B(b[27]), .Z(N34) );
  XOR2_X1 U1165 ( .A(n197), .B(b[28]), .Z(N33) );
  XOR2_X1 U1166 ( .A(n197), .B(b[29]), .Z(N32) );
  XOR2_X1 U1167 ( .A(n197), .B(b[30]), .Z(N31) );
  XOR2_X1 U1168 ( .A(a[31]), .B(a[0]), .Z(N30) );
  XOR2_X1 U1169 ( .A(n4), .B(a[27]), .Z(N3) );
  XOR2_X1 U1171 ( .A(n5), .B(a[2]), .Z(N28) );
  XOR2_X1 U1172 ( .A(a[3]), .B(n7), .Z(N27) );
  XOR2_X1 U1173 ( .A(a[4]), .B(n6), .Z(N26) );
  XOR2_X1 U1174 ( .A(a[5]), .B(n7), .Z(N25) );
  XOR2_X1 U1175 ( .A(a[6]), .B(n6), .Z(N24) );
  XOR2_X1 U1176 ( .A(a[7]), .B(n7), .Z(N23) );
  XOR2_X1 U1177 ( .A(a[8]), .B(n6), .Z(N22) );
  XOR2_X1 U1178 ( .A(a[9]), .B(n7), .Z(N21) );
  XOR2_X1 U1179 ( .A(n4), .B(a[10]), .Z(N20) );
  XOR2_X1 U1180 ( .A(n5), .B(a[28]), .Z(N2) );
  XOR2_X1 U1181 ( .A(n5), .B(a[11]), .Z(N19) );
  XOR2_X1 U1182 ( .A(n4), .B(a[12]), .Z(N18) );
  XOR2_X1 U1183 ( .A(n5), .B(a[13]), .Z(N17) );
  XOR2_X1 U1184 ( .A(n4), .B(a[14]), .Z(N16) );
  XOR2_X1 U1185 ( .A(n6), .B(a[15]), .Z(N15) );
  XOR2_X1 U1186 ( .A(n7), .B(a[16]), .Z(N14) );
  XOR2_X1 U1187 ( .A(n6), .B(a[17]), .Z(N13) );
  XOR2_X1 U1188 ( .A(n68), .B(n195), .Z(N125) );
  XOR2_X1 U1189 ( .A(tempResult[1]), .B(n195), .Z(N124) );
  XOR2_X1 U1190 ( .A(tempResult[2]), .B(n195), .Z(N123) );
  XOR2_X1 U1191 ( .A(tempResult[3]), .B(n195), .Z(N122) );
  XOR2_X1 U1192 ( .A(tempResult[4]), .B(n195), .Z(N121) );
  XOR2_X1 U1193 ( .A(tempResult[5]), .B(n195), .Z(N120) );
  XOR2_X1 U1194 ( .A(n7), .B(a[18]), .Z(N12) );
  XOR2_X1 U1195 ( .A(tempResult[6]), .B(n195), .Z(N119) );
  XOR2_X1 U1196 ( .A(tempResult[7]), .B(n195), .Z(N118) );
  XOR2_X1 U1197 ( .A(tempResult[8]), .B(n195), .Z(N117) );
  XOR2_X1 U1198 ( .A(tempResult[9]), .B(n195), .Z(N116) );
  XOR2_X1 U1199 ( .A(tempResult[10]), .B(n195), .Z(N115) );
  XOR2_X1 U1200 ( .A(tempResult[11]), .B(n195), .Z(N114) );
  XOR2_X1 U1201 ( .A(tempResult[12]), .B(n196), .Z(N113) );
  XOR2_X1 U1202 ( .A(tempResult[13]), .B(n196), .Z(N112) );
  XOR2_X1 U1203 ( .A(tempResult[14]), .B(n196), .Z(N111) );
  XOR2_X1 U1204 ( .A(tempResult[15]), .B(n196), .Z(N110) );
  XOR2_X1 U1205 ( .A(n6), .B(a[19]), .Z(N11) );
  XOR2_X1 U1206 ( .A(tempResult[16]), .B(n196), .Z(N109) );
  XOR2_X1 U1207 ( .A(tempResult[17]), .B(n196), .Z(N108) );
  XOR2_X1 U1208 ( .A(tempResult[18]), .B(n196), .Z(N107) );
  XOR2_X1 U1209 ( .A(tempResult[19]), .B(n196), .Z(N106) );
  XOR2_X1 U1210 ( .A(tempResult[20]), .B(n196), .Z(N105) );
  XOR2_X1 U1211 ( .A(tempResult[21]), .B(n196), .Z(N104) );
  XOR2_X1 U1212 ( .A(tempResult[22]), .B(n196), .Z(N103) );
  XOR2_X1 U1213 ( .A(tempResult[23]), .B(n196), .Z(N102) );
  XOR2_X1 U1214 ( .A(tempResult[24]), .B(n196), .Z(N101) );
  XOR2_X1 U1215 ( .A(tempResult[25]), .B(n196), .Z(N100) );
  XOR2_X1 U1216 ( .A(n6), .B(n197), .Z(finalSign) );
  XOR2_X1 U1217 ( .A(n7), .B(a[20]), .Z(N10) );
  XOR2_X1 U1218 ( .A(n7), .B(a[29]), .Z(N1) );
  XOR2_X1 U1219 ( .A(n4), .B(a[30]), .Z(N0) );
  carryLookAheadAdder_0 A0 ( .a({1'b0, tempResultA_0__30_, tempResultA_0__29_, 
        tempResultA_0__28_, tempResultA_0__27_, tempResultA_0__26_, 
        tempResultA_0__25_, tempResultA_0__24_, tempResultA_0__23_, 
        tempResultA_0__22_, tempResultA_0__21_, tempResultA_0__20_, 
        tempResultA_0__19_, tempResultA_0__18_, tempResultA_0__17_, 
        tempResultA_0__16_, tempResultA_0__15_, tempResultA_0__14_, 
        tempResultA_0__13_, tempResultA_0__12_, tempResultA_0__11_, 
        tempResultA_0__10_, tempResultA_0__9_, tempResultA_0__8_, 
        tempResultA_0__7_, tempResultA_0__6_, tempResultA_0__5_, 
        tempResultA_0__4_, tempResultA_0__3_, tempResultA_0__2_, 
        tempResultA_0__1_, tempResultA_0__0_}), .b(tempResultB[31:0]), .cin(
        1'b0), .result({tempResultA_1__30_, tempResultA_1__29_, 
        tempResultA_1__28_, tempResultA_1__27_, tempResultA_1__26_, 
        tempResultA_1__25_, tempResultA_1__24_, tempResultA_1__23_, 
        tempResultA_1__22_, tempResultA_1__21_, tempResultA_1__20_, 
        tempResultA_1__19_, tempResultA_1__18_, tempResultA_1__17_, 
        tempResultA_1__16_, tempResultA_1__15_, tempResultA_1__14_, 
        tempResultA_1__13_, tempResultA_1__12_, tempResultA_1__11_, 
        tempResultA_1__10_, tempResultA_1__9_, tempResultA_1__8_, 
        tempResultA_1__7_, tempResultA_1__6_, tempResultA_1__5_, 
        tempResultA_1__4_, tempResultA_1__3_, tempResultA_1__2_, 
        tempResultA_1__1_, tempResultA_1__0_, tempResult[1]}), .cout(
        tempResultA_1__31_) );
  carryLookAheadAdder_30 generating_partialProducts_1__A1 ( .a({
        tempResultA_1__31_, tempResultA_1__30_, tempResultA_1__29_, 
        tempResultA_1__28_, tempResultA_1__27_, tempResultA_1__26_, 
        tempResultA_1__25_, tempResultA_1__24_, tempResultA_1__23_, 
        tempResultA_1__22_, tempResultA_1__21_, tempResultA_1__20_, 
        tempResultA_1__19_, tempResultA_1__18_, tempResultA_1__17_, 
        tempResultA_1__16_, tempResultA_1__15_, tempResultA_1__14_, 
        tempResultA_1__13_, tempResultA_1__12_, tempResultA_1__11_, 
        tempResultA_1__10_, tempResultA_1__9_, tempResultA_1__8_, 
        tempResultA_1__7_, tempResultA_1__6_, tempResultA_1__5_, 
        tempResultA_1__4_, tempResultA_1__3_, tempResultA_1__2_, 
        tempResultA_1__1_, tempResultA_1__0_}), .b(tempResultB[63:32]), .cin(
        1'b0), .result({tempResultA_2__30_, tempResultA_2__29_, 
        tempResultA_2__28_, tempResultA_2__27_, tempResultA_2__26_, 
        tempResultA_2__25_, tempResultA_2__24_, tempResultA_2__23_, 
        tempResultA_2__22_, tempResultA_2__21_, tempResultA_2__20_, 
        tempResultA_2__19_, tempResultA_2__18_, tempResultA_2__17_, 
        tempResultA_2__16_, tempResultA_2__15_, tempResultA_2__14_, 
        tempResultA_2__13_, tempResultA_2__12_, tempResultA_2__11_, 
        tempResultA_2__10_, tempResultA_2__9_, tempResultA_2__8_, 
        tempResultA_2__7_, tempResultA_2__6_, tempResultA_2__5_, 
        tempResultA_2__4_, tempResultA_2__3_, tempResultA_2__2_, 
        tempResultA_2__1_, tempResultA_2__0_, tempResult[2]}), .cout(
        tempResultA_2__31_) );
  carryLookAheadAdder_29 generating_partialProducts_2__A1 ( .a({
        tempResultA_2__31_, tempResultA_2__30_, tempResultA_2__29_, 
        tempResultA_2__28_, tempResultA_2__27_, tempResultA_2__26_, 
        tempResultA_2__25_, tempResultA_2__24_, tempResultA_2__23_, 
        tempResultA_2__22_, tempResultA_2__21_, tempResultA_2__20_, 
        tempResultA_2__19_, tempResultA_2__18_, tempResultA_2__17_, 
        tempResultA_2__16_, tempResultA_2__15_, tempResultA_2__14_, 
        tempResultA_2__13_, tempResultA_2__12_, tempResultA_2__11_, 
        tempResultA_2__10_, tempResultA_2__9_, tempResultA_2__8_, 
        tempResultA_2__7_, tempResultA_2__6_, tempResultA_2__5_, 
        tempResultA_2__4_, tempResultA_2__3_, tempResultA_2__2_, 
        tempResultA_2__1_, tempResultA_2__0_}), .b(tempResultB[95:64]), .cin(
        1'b0), .result({tempResultA_3__30_, tempResultA_3__29_, 
        tempResultA_3__28_, tempResultA_3__27_, tempResultA_3__26_, 
        tempResultA_3__25_, tempResultA_3__24_, tempResultA_3__23_, 
        tempResultA_3__22_, tempResultA_3__21_, tempResultA_3__20_, 
        tempResultA_3__19_, tempResultA_3__18_, tempResultA_3__17_, 
        tempResultA_3__16_, tempResultA_3__15_, tempResultA_3__14_, 
        tempResultA_3__13_, tempResultA_3__12_, tempResultA_3__11_, 
        tempResultA_3__10_, tempResultA_3__9_, tempResultA_3__8_, 
        tempResultA_3__7_, tempResultA_3__6_, tempResultA_3__5_, 
        tempResultA_3__4_, tempResultA_3__3_, tempResultA_3__2_, 
        tempResultA_3__1_, tempResultA_3__0_, tempResult[3]}), .cout(
        tempResultA_3__31_) );
  carryLookAheadAdder_28 generating_partialProducts_3__A1 ( .a({
        tempResultA_3__31_, tempResultA_3__30_, tempResultA_3__29_, 
        tempResultA_3__28_, tempResultA_3__27_, tempResultA_3__26_, 
        tempResultA_3__25_, tempResultA_3__24_, tempResultA_3__23_, 
        tempResultA_3__22_, tempResultA_3__21_, tempResultA_3__20_, 
        tempResultA_3__19_, tempResultA_3__18_, tempResultA_3__17_, 
        tempResultA_3__16_, tempResultA_3__15_, tempResultA_3__14_, 
        tempResultA_3__13_, tempResultA_3__12_, tempResultA_3__11_, 
        tempResultA_3__10_, tempResultA_3__9_, tempResultA_3__8_, 
        tempResultA_3__7_, tempResultA_3__6_, tempResultA_3__5_, 
        tempResultA_3__4_, tempResultA_3__3_, tempResultA_3__2_, 
        tempResultA_3__1_, tempResultA_3__0_}), .b(tempResultB[127:96]), .cin(
        1'b0), .result({tempResultA_4__30_, tempResultA_4__29_, 
        tempResultA_4__28_, tempResultA_4__27_, tempResultA_4__26_, 
        tempResultA_4__25_, tempResultA_4__24_, tempResultA_4__23_, 
        tempResultA_4__22_, tempResultA_4__21_, tempResultA_4__20_, 
        tempResultA_4__19_, tempResultA_4__18_, tempResultA_4__17_, 
        tempResultA_4__16_, tempResultA_4__15_, tempResultA_4__14_, 
        tempResultA_4__13_, tempResultA_4__12_, tempResultA_4__11_, 
        tempResultA_4__10_, tempResultA_4__9_, tempResultA_4__8_, 
        tempResultA_4__7_, tempResultA_4__6_, tempResultA_4__5_, 
        tempResultA_4__4_, tempResultA_4__3_, tempResultA_4__2_, 
        tempResultA_4__1_, tempResultA_4__0_, tempResult[4]}), .cout(
        tempResultA_4__31_) );
  carryLookAheadAdder_27 generating_partialProducts_4__A1 ( .a({
        tempResultA_4__31_, tempResultA_4__30_, tempResultA_4__29_, 
        tempResultA_4__28_, tempResultA_4__27_, tempResultA_4__26_, 
        tempResultA_4__25_, tempResultA_4__24_, tempResultA_4__23_, 
        tempResultA_4__22_, tempResultA_4__21_, tempResultA_4__20_, 
        tempResultA_4__19_, tempResultA_4__18_, tempResultA_4__17_, 
        tempResultA_4__16_, tempResultA_4__15_, tempResultA_4__14_, 
        tempResultA_4__13_, tempResultA_4__12_, tempResultA_4__11_, 
        tempResultA_4__10_, tempResultA_4__9_, tempResultA_4__8_, 
        tempResultA_4__7_, tempResultA_4__6_, tempResultA_4__5_, 
        tempResultA_4__4_, tempResultA_4__3_, tempResultA_4__2_, 
        tempResultA_4__1_, tempResultA_4__0_}), .b(tempResultB[159:128]), 
        .cin(1'b0), .result({tempResultA_5__30_, tempResultA_5__29_, 
        tempResultA_5__28_, tempResultA_5__27_, tempResultA_5__26_, 
        tempResultA_5__25_, tempResultA_5__24_, tempResultA_5__23_, 
        tempResultA_5__22_, tempResultA_5__21_, tempResultA_5__20_, 
        tempResultA_5__19_, tempResultA_5__18_, tempResultA_5__17_, 
        tempResultA_5__16_, tempResultA_5__15_, tempResultA_5__14_, 
        tempResultA_5__13_, tempResultA_5__12_, tempResultA_5__11_, 
        tempResultA_5__10_, tempResultA_5__9_, tempResultA_5__8_, 
        tempResultA_5__7_, tempResultA_5__6_, tempResultA_5__5_, 
        tempResultA_5__4_, tempResultA_5__3_, tempResultA_5__2_, 
        tempResultA_5__1_, tempResultA_5__0_, tempResult[5]}), .cout(
        tempResultA_5__31_) );
  carryLookAheadAdder_26 generating_partialProducts_5__A1 ( .a({
        tempResultA_5__31_, tempResultA_5__30_, tempResultA_5__29_, 
        tempResultA_5__28_, tempResultA_5__27_, tempResultA_5__26_, 
        tempResultA_5__25_, tempResultA_5__24_, tempResultA_5__23_, 
        tempResultA_5__22_, tempResultA_5__21_, tempResultA_5__20_, 
        tempResultA_5__19_, tempResultA_5__18_, tempResultA_5__17_, 
        tempResultA_5__16_, tempResultA_5__15_, tempResultA_5__14_, 
        tempResultA_5__13_, tempResultA_5__12_, tempResultA_5__11_, 
        tempResultA_5__10_, tempResultA_5__9_, tempResultA_5__8_, 
        tempResultA_5__7_, tempResultA_5__6_, tempResultA_5__5_, 
        tempResultA_5__4_, tempResultA_5__3_, tempResultA_5__2_, 
        tempResultA_5__1_, tempResultA_5__0_}), .b(tempResultB[191:160]), 
        .cin(1'b0), .result({tempResultA_6__30_, tempResultA_6__29_, 
        tempResultA_6__28_, tempResultA_6__27_, tempResultA_6__26_, 
        tempResultA_6__25_, tempResultA_6__24_, tempResultA_6__23_, 
        tempResultA_6__22_, tempResultA_6__21_, tempResultA_6__20_, 
        tempResultA_6__19_, tempResultA_6__18_, tempResultA_6__17_, 
        tempResultA_6__16_, tempResultA_6__15_, tempResultA_6__14_, 
        tempResultA_6__13_, tempResultA_6__12_, tempResultA_6__11_, 
        tempResultA_6__10_, tempResultA_6__9_, tempResultA_6__8_, 
        tempResultA_6__7_, tempResultA_6__6_, tempResultA_6__5_, 
        tempResultA_6__4_, tempResultA_6__3_, tempResultA_6__2_, 
        tempResultA_6__1_, tempResultA_6__0_, tempResult[6]}), .cout(
        tempResultA_6__31_) );
  carryLookAheadAdder_25 generating_partialProducts_6__A1 ( .a({
        tempResultA_6__31_, tempResultA_6__30_, tempResultA_6__29_, 
        tempResultA_6__28_, tempResultA_6__27_, tempResultA_6__26_, 
        tempResultA_6__25_, tempResultA_6__24_, tempResultA_6__23_, 
        tempResultA_6__22_, tempResultA_6__21_, tempResultA_6__20_, 
        tempResultA_6__19_, tempResultA_6__18_, tempResultA_6__17_, 
        tempResultA_6__16_, tempResultA_6__15_, tempResultA_6__14_, 
        tempResultA_6__13_, tempResultA_6__12_, tempResultA_6__11_, 
        tempResultA_6__10_, tempResultA_6__9_, tempResultA_6__8_, 
        tempResultA_6__7_, tempResultA_6__6_, tempResultA_6__5_, 
        tempResultA_6__4_, tempResultA_6__3_, tempResultA_6__2_, 
        tempResultA_6__1_, tempResultA_6__0_}), .b(tempResultB[223:192]), 
        .cin(1'b0), .result({tempResultA_7__30_, tempResultA_7__29_, 
        tempResultA_7__28_, tempResultA_7__27_, tempResultA_7__26_, 
        tempResultA_7__25_, tempResultA_7__24_, tempResultA_7__23_, 
        tempResultA_7__22_, tempResultA_7__21_, tempResultA_7__20_, 
        tempResultA_7__19_, tempResultA_7__18_, tempResultA_7__17_, 
        tempResultA_7__16_, tempResultA_7__15_, tempResultA_7__14_, 
        tempResultA_7__13_, tempResultA_7__12_, tempResultA_7__11_, 
        tempResultA_7__10_, tempResultA_7__9_, tempResultA_7__8_, 
        tempResultA_7__7_, tempResultA_7__6_, tempResultA_7__5_, 
        tempResultA_7__4_, tempResultA_7__3_, tempResultA_7__2_, 
        tempResultA_7__1_, tempResultA_7__0_, tempResult[7]}), .cout(
        tempResultA_7__31_) );
  carryLookAheadAdder_24 generating_partialProducts_7__A1 ( .a({
        tempResultA_7__31_, tempResultA_7__30_, tempResultA_7__29_, 
        tempResultA_7__28_, tempResultA_7__27_, tempResultA_7__26_, 
        tempResultA_7__25_, tempResultA_7__24_, tempResultA_7__23_, 
        tempResultA_7__22_, tempResultA_7__21_, tempResultA_7__20_, 
        tempResultA_7__19_, tempResultA_7__18_, tempResultA_7__17_, 
        tempResultA_7__16_, tempResultA_7__15_, tempResultA_7__14_, 
        tempResultA_7__13_, tempResultA_7__12_, tempResultA_7__11_, 
        tempResultA_7__10_, tempResultA_7__9_, tempResultA_7__8_, 
        tempResultA_7__7_, tempResultA_7__6_, tempResultA_7__5_, 
        tempResultA_7__4_, tempResultA_7__3_, tempResultA_7__2_, 
        tempResultA_7__1_, tempResultA_7__0_}), .b(tempResultB[255:224]), 
        .cin(1'b0), .result({tempResultA_8__30_, tempResultA_8__29_, 
        tempResultA_8__28_, tempResultA_8__27_, tempResultA_8__26_, 
        tempResultA_8__25_, tempResultA_8__24_, tempResultA_8__23_, 
        tempResultA_8__22_, tempResultA_8__21_, tempResultA_8__20_, 
        tempResultA_8__19_, tempResultA_8__18_, tempResultA_8__17_, 
        tempResultA_8__16_, tempResultA_8__15_, tempResultA_8__14_, 
        tempResultA_8__13_, tempResultA_8__12_, tempResultA_8__11_, 
        tempResultA_8__10_, tempResultA_8__9_, tempResultA_8__8_, 
        tempResultA_8__7_, tempResultA_8__6_, tempResultA_8__5_, 
        tempResultA_8__4_, tempResultA_8__3_, tempResultA_8__2_, 
        tempResultA_8__1_, tempResultA_8__0_, tempResult[8]}), .cout(
        tempResultA_8__31_) );
  carryLookAheadAdder_23 generating_partialProducts_8__A1 ( .a({
        tempResultA_8__31_, tempResultA_8__30_, tempResultA_8__29_, 
        tempResultA_8__28_, tempResultA_8__27_, tempResultA_8__26_, 
        tempResultA_8__25_, tempResultA_8__24_, tempResultA_8__23_, 
        tempResultA_8__22_, tempResultA_8__21_, tempResultA_8__20_, 
        tempResultA_8__19_, tempResultA_8__18_, tempResultA_8__17_, 
        tempResultA_8__16_, tempResultA_8__15_, tempResultA_8__14_, 
        tempResultA_8__13_, tempResultA_8__12_, tempResultA_8__11_, 
        tempResultA_8__10_, tempResultA_8__9_, tempResultA_8__8_, 
        tempResultA_8__7_, tempResultA_8__6_, tempResultA_8__5_, 
        tempResultA_8__4_, tempResultA_8__3_, tempResultA_8__2_, 
        tempResultA_8__1_, tempResultA_8__0_}), .b(tempResultB[287:256]), 
        .cin(1'b0), .result({tempResultA_9__30_, tempResultA_9__29_, 
        tempResultA_9__28_, tempResultA_9__27_, tempResultA_9__26_, 
        tempResultA_9__25_, tempResultA_9__24_, tempResultA_9__23_, 
        tempResultA_9__22_, tempResultA_9__21_, tempResultA_9__20_, 
        tempResultA_9__19_, tempResultA_9__18_, tempResultA_9__17_, 
        tempResultA_9__16_, tempResultA_9__15_, tempResultA_9__14_, 
        tempResultA_9__13_, tempResultA_9__12_, tempResultA_9__11_, 
        tempResultA_9__10_, tempResultA_9__9_, tempResultA_9__8_, 
        tempResultA_9__7_, tempResultA_9__6_, tempResultA_9__5_, 
        tempResultA_9__4_, tempResultA_9__3_, tempResultA_9__2_, 
        tempResultA_9__1_, tempResultA_9__0_, tempResult[9]}), .cout(
        tempResultA_9__31_) );
  carryLookAheadAdder_22 generating_partialProducts_9__A1 ( .a({
        tempResultA_9__31_, tempResultA_9__30_, tempResultA_9__29_, 
        tempResultA_9__28_, tempResultA_9__27_, tempResultA_9__26_, 
        tempResultA_9__25_, tempResultA_9__24_, tempResultA_9__23_, 
        tempResultA_9__22_, tempResultA_9__21_, tempResultA_9__20_, 
        tempResultA_9__19_, tempResultA_9__18_, tempResultA_9__17_, 
        tempResultA_9__16_, tempResultA_9__15_, tempResultA_9__14_, 
        tempResultA_9__13_, tempResultA_9__12_, tempResultA_9__11_, 
        tempResultA_9__10_, tempResultA_9__9_, tempResultA_9__8_, 
        tempResultA_9__7_, tempResultA_9__6_, tempResultA_9__5_, 
        tempResultA_9__4_, tempResultA_9__3_, tempResultA_9__2_, 
        tempResultA_9__1_, tempResultA_9__0_}), .b(tempResultB[319:288]), 
        .cin(1'b0), .result({tempResultA_10__30_, tempResultA_10__29_, 
        tempResultA_10__28_, tempResultA_10__27_, tempResultA_10__26_, 
        tempResultA_10__25_, tempResultA_10__24_, tempResultA_10__23_, 
        tempResultA_10__22_, tempResultA_10__21_, tempResultA_10__20_, 
        tempResultA_10__19_, tempResultA_10__18_, tempResultA_10__17_, 
        tempResultA_10__16_, tempResultA_10__15_, tempResultA_10__14_, 
        tempResultA_10__13_, tempResultA_10__12_, tempResultA_10__11_, 
        tempResultA_10__10_, tempResultA_10__9_, tempResultA_10__8_, 
        tempResultA_10__7_, tempResultA_10__6_, tempResultA_10__5_, 
        tempResultA_10__4_, tempResultA_10__3_, tempResultA_10__2_, 
        tempResultA_10__1_, tempResultA_10__0_, tempResult[10]}), .cout(
        tempResultA_10__31_) );
  carryLookAheadAdder_21 generating_partialProducts_10__A1 ( .a({
        tempResultA_10__31_, tempResultA_10__30_, tempResultA_10__29_, 
        tempResultA_10__28_, tempResultA_10__27_, tempResultA_10__26_, 
        tempResultA_10__25_, tempResultA_10__24_, tempResultA_10__23_, 
        tempResultA_10__22_, tempResultA_10__21_, tempResultA_10__20_, 
        tempResultA_10__19_, tempResultA_10__18_, tempResultA_10__17_, 
        tempResultA_10__16_, tempResultA_10__15_, tempResultA_10__14_, 
        tempResultA_10__13_, tempResultA_10__12_, tempResultA_10__11_, 
        tempResultA_10__10_, tempResultA_10__9_, tempResultA_10__8_, 
        tempResultA_10__7_, tempResultA_10__6_, tempResultA_10__5_, 
        tempResultA_10__4_, tempResultA_10__3_, tempResultA_10__2_, 
        tempResultA_10__1_, tempResultA_10__0_}), .b(tempResultB[351:320]), 
        .cin(1'b0), .result({tempResultA_11__30_, tempResultA_11__29_, 
        tempResultA_11__28_, tempResultA_11__27_, tempResultA_11__26_, 
        tempResultA_11__25_, tempResultA_11__24_, tempResultA_11__23_, 
        tempResultA_11__22_, tempResultA_11__21_, tempResultA_11__20_, 
        tempResultA_11__19_, tempResultA_11__18_, tempResultA_11__17_, 
        tempResultA_11__16_, tempResultA_11__15_, tempResultA_11__14_, 
        tempResultA_11__13_, tempResultA_11__12_, tempResultA_11__11_, 
        tempResultA_11__10_, tempResultA_11__9_, tempResultA_11__8_, 
        tempResultA_11__7_, tempResultA_11__6_, tempResultA_11__5_, 
        tempResultA_11__4_, tempResultA_11__3_, tempResultA_11__2_, 
        tempResultA_11__1_, tempResultA_11__0_, tempResult[11]}), .cout(
        tempResultA_11__31_) );
  carryLookAheadAdder_20 generating_partialProducts_11__A1 ( .a({
        tempResultA_11__31_, tempResultA_11__30_, tempResultA_11__29_, 
        tempResultA_11__28_, tempResultA_11__27_, tempResultA_11__26_, 
        tempResultA_11__25_, tempResultA_11__24_, tempResultA_11__23_, 
        tempResultA_11__22_, tempResultA_11__21_, tempResultA_11__20_, 
        tempResultA_11__19_, tempResultA_11__18_, tempResultA_11__17_, 
        tempResultA_11__16_, tempResultA_11__15_, tempResultA_11__14_, 
        tempResultA_11__13_, tempResultA_11__12_, tempResultA_11__11_, 
        tempResultA_11__10_, tempResultA_11__9_, tempResultA_11__8_, 
        tempResultA_11__7_, tempResultA_11__6_, tempResultA_11__5_, 
        tempResultA_11__4_, tempResultA_11__3_, tempResultA_11__2_, 
        tempResultA_11__1_, tempResultA_11__0_}), .b(tempResultB[383:352]), 
        .cin(1'b0), .result({tempResultA_12__30_, tempResultA_12__29_, 
        tempResultA_12__28_, tempResultA_12__27_, tempResultA_12__26_, 
        tempResultA_12__25_, tempResultA_12__24_, tempResultA_12__23_, 
        tempResultA_12__22_, tempResultA_12__21_, tempResultA_12__20_, 
        tempResultA_12__19_, tempResultA_12__18_, tempResultA_12__17_, 
        tempResultA_12__16_, tempResultA_12__15_, tempResultA_12__14_, 
        tempResultA_12__13_, tempResultA_12__12_, tempResultA_12__11_, 
        tempResultA_12__10_, tempResultA_12__9_, tempResultA_12__8_, 
        tempResultA_12__7_, tempResultA_12__6_, tempResultA_12__5_, 
        tempResultA_12__4_, tempResultA_12__3_, tempResultA_12__2_, 
        tempResultA_12__1_, tempResultA_12__0_, tempResult[12]}), .cout(
        tempResultA_12__31_) );
  carryLookAheadAdder_19 generating_partialProducts_12__A1 ( .a({
        tempResultA_12__31_, tempResultA_12__30_, tempResultA_12__29_, 
        tempResultA_12__28_, tempResultA_12__27_, tempResultA_12__26_, 
        tempResultA_12__25_, tempResultA_12__24_, tempResultA_12__23_, 
        tempResultA_12__22_, tempResultA_12__21_, tempResultA_12__20_, 
        tempResultA_12__19_, tempResultA_12__18_, tempResultA_12__17_, 
        tempResultA_12__16_, tempResultA_12__15_, tempResultA_12__14_, 
        tempResultA_12__13_, tempResultA_12__12_, tempResultA_12__11_, 
        tempResultA_12__10_, tempResultA_12__9_, tempResultA_12__8_, 
        tempResultA_12__7_, tempResultA_12__6_, tempResultA_12__5_, 
        tempResultA_12__4_, tempResultA_12__3_, tempResultA_12__2_, 
        tempResultA_12__1_, tempResultA_12__0_}), .b(tempResultB[415:384]), 
        .cin(1'b0), .result({tempResultA_13__30_, tempResultA_13__29_, 
        tempResultA_13__28_, tempResultA_13__27_, tempResultA_13__26_, 
        tempResultA_13__25_, tempResultA_13__24_, tempResultA_13__23_, 
        tempResultA_13__22_, tempResultA_13__21_, tempResultA_13__20_, 
        tempResultA_13__19_, tempResultA_13__18_, tempResultA_13__17_, 
        tempResultA_13__16_, tempResultA_13__15_, tempResultA_13__14_, 
        tempResultA_13__13_, tempResultA_13__12_, tempResultA_13__11_, 
        tempResultA_13__10_, tempResultA_13__9_, tempResultA_13__8_, 
        tempResultA_13__7_, tempResultA_13__6_, tempResultA_13__5_, 
        tempResultA_13__4_, tempResultA_13__3_, tempResultA_13__2_, 
        tempResultA_13__1_, tempResultA_13__0_, tempResult[13]}), .cout(
        tempResultA_13__31_) );
  carryLookAheadAdder_18 generating_partialProducts_13__A1 ( .a({
        tempResultA_13__31_, tempResultA_13__30_, tempResultA_13__29_, 
        tempResultA_13__28_, tempResultA_13__27_, tempResultA_13__26_, 
        tempResultA_13__25_, tempResultA_13__24_, tempResultA_13__23_, 
        tempResultA_13__22_, tempResultA_13__21_, tempResultA_13__20_, 
        tempResultA_13__19_, tempResultA_13__18_, tempResultA_13__17_, 
        tempResultA_13__16_, tempResultA_13__15_, tempResultA_13__14_, 
        tempResultA_13__13_, tempResultA_13__12_, tempResultA_13__11_, 
        tempResultA_13__10_, tempResultA_13__9_, tempResultA_13__8_, 
        tempResultA_13__7_, tempResultA_13__6_, tempResultA_13__5_, 
        tempResultA_13__4_, tempResultA_13__3_, tempResultA_13__2_, 
        tempResultA_13__1_, tempResultA_13__0_}), .b(tempResultB[447:416]), 
        .cin(1'b0), .result({tempResultA_14__30_, tempResultA_14__29_, 
        tempResultA_14__28_, tempResultA_14__27_, tempResultA_14__26_, 
        tempResultA_14__25_, tempResultA_14__24_, tempResultA_14__23_, 
        tempResultA_14__22_, tempResultA_14__21_, tempResultA_14__20_, 
        tempResultA_14__19_, tempResultA_14__18_, tempResultA_14__17_, 
        tempResultA_14__16_, tempResultA_14__15_, tempResultA_14__14_, 
        tempResultA_14__13_, tempResultA_14__12_, tempResultA_14__11_, 
        tempResultA_14__10_, tempResultA_14__9_, tempResultA_14__8_, 
        tempResultA_14__7_, tempResultA_14__6_, tempResultA_14__5_, 
        tempResultA_14__4_, tempResultA_14__3_, tempResultA_14__2_, 
        tempResultA_14__1_, tempResultA_14__0_, tempResult[14]}), .cout(
        tempResultA_14__31_) );
  carryLookAheadAdder_17 generating_partialProducts_14__A1 ( .a({
        tempResultA_14__31_, tempResultA_14__30_, tempResultA_14__29_, 
        tempResultA_14__28_, tempResultA_14__27_, tempResultA_14__26_, 
        tempResultA_14__25_, tempResultA_14__24_, tempResultA_14__23_, 
        tempResultA_14__22_, tempResultA_14__21_, tempResultA_14__20_, 
        tempResultA_14__19_, tempResultA_14__18_, tempResultA_14__17_, 
        tempResultA_14__16_, tempResultA_14__15_, tempResultA_14__14_, 
        tempResultA_14__13_, tempResultA_14__12_, tempResultA_14__11_, 
        tempResultA_14__10_, tempResultA_14__9_, tempResultA_14__8_, 
        tempResultA_14__7_, tempResultA_14__6_, tempResultA_14__5_, 
        tempResultA_14__4_, tempResultA_14__3_, tempResultA_14__2_, 
        tempResultA_14__1_, tempResultA_14__0_}), .b(tempResultB[479:448]), 
        .cin(1'b0), .result({tempResultA_15__30_, tempResultA_15__29_, 
        tempResultA_15__28_, tempResultA_15__27_, tempResultA_15__26_, 
        tempResultA_15__25_, tempResultA_15__24_, tempResultA_15__23_, 
        tempResultA_15__22_, tempResultA_15__21_, tempResultA_15__20_, 
        tempResultA_15__19_, tempResultA_15__18_, tempResultA_15__17_, 
        tempResultA_15__16_, tempResultA_15__15_, tempResultA_15__14_, 
        tempResultA_15__13_, tempResultA_15__12_, tempResultA_15__11_, 
        tempResultA_15__10_, tempResultA_15__9_, tempResultA_15__8_, 
        tempResultA_15__7_, tempResultA_15__6_, tempResultA_15__5_, 
        tempResultA_15__4_, tempResultA_15__3_, tempResultA_15__2_, 
        tempResultA_15__1_, tempResultA_15__0_, tempResult[15]}), .cout(
        tempResultA_15__31_) );
  carryLookAheadAdder_16 generating_partialProducts_15__A1 ( .a({
        tempResultA_15__31_, tempResultA_15__30_, tempResultA_15__29_, 
        tempResultA_15__28_, tempResultA_15__27_, tempResultA_15__26_, 
        tempResultA_15__25_, tempResultA_15__24_, tempResultA_15__23_, 
        tempResultA_15__22_, tempResultA_15__21_, tempResultA_15__20_, 
        tempResultA_15__19_, tempResultA_15__18_, tempResultA_15__17_, 
        tempResultA_15__16_, tempResultA_15__15_, tempResultA_15__14_, 
        tempResultA_15__13_, tempResultA_15__12_, tempResultA_15__11_, 
        tempResultA_15__10_, tempResultA_15__9_, tempResultA_15__8_, 
        tempResultA_15__7_, tempResultA_15__6_, tempResultA_15__5_, 
        tempResultA_15__4_, tempResultA_15__3_, tempResultA_15__2_, 
        tempResultA_15__1_, tempResultA_15__0_}), .b(tempResultB[511:480]), 
        .cin(1'b0), .result({tempResultA_16__30_, tempResultA_16__29_, 
        tempResultA_16__28_, tempResultA_16__27_, tempResultA_16__26_, 
        tempResultA_16__25_, tempResultA_16__24_, tempResultA_16__23_, 
        tempResultA_16__22_, tempResultA_16__21_, tempResultA_16__20_, 
        tempResultA_16__19_, tempResultA_16__18_, tempResultA_16__17_, 
        tempResultA_16__16_, tempResultA_16__15_, tempResultA_16__14_, 
        tempResultA_16__13_, tempResultA_16__12_, tempResultA_16__11_, 
        tempResultA_16__10_, tempResultA_16__9_, tempResultA_16__8_, 
        tempResultA_16__7_, tempResultA_16__6_, tempResultA_16__5_, 
        tempResultA_16__4_, tempResultA_16__3_, tempResultA_16__2_, 
        tempResultA_16__1_, tempResultA_16__0_, tempResult[16]}), .cout(
        tempResultA_16__31_) );
  carryLookAheadAdder_15 generating_partialProducts_16__A1 ( .a({
        tempResultA_16__31_, tempResultA_16__30_, tempResultA_16__29_, 
        tempResultA_16__28_, tempResultA_16__27_, tempResultA_16__26_, 
        tempResultA_16__25_, tempResultA_16__24_, tempResultA_16__23_, 
        tempResultA_16__22_, tempResultA_16__21_, tempResultA_16__20_, 
        tempResultA_16__19_, tempResultA_16__18_, tempResultA_16__17_, 
        tempResultA_16__16_, tempResultA_16__15_, tempResultA_16__14_, 
        tempResultA_16__13_, tempResultA_16__12_, tempResultA_16__11_, 
        tempResultA_16__10_, tempResultA_16__9_, tempResultA_16__8_, 
        tempResultA_16__7_, tempResultA_16__6_, tempResultA_16__5_, 
        tempResultA_16__4_, tempResultA_16__3_, tempResultA_16__2_, 
        tempResultA_16__1_, tempResultA_16__0_}), .b(tempResultB[543:512]), 
        .cin(1'b0), .result({tempResultA_17__30_, tempResultA_17__29_, 
        tempResultA_17__28_, tempResultA_17__27_, tempResultA_17__26_, 
        tempResultA_17__25_, tempResultA_17__24_, tempResultA_17__23_, 
        tempResultA_17__22_, tempResultA_17__21_, tempResultA_17__20_, 
        tempResultA_17__19_, tempResultA_17__18_, tempResultA_17__17_, 
        tempResultA_17__16_, tempResultA_17__15_, tempResultA_17__14_, 
        tempResultA_17__13_, tempResultA_17__12_, tempResultA_17__11_, 
        tempResultA_17__10_, tempResultA_17__9_, tempResultA_17__8_, 
        tempResultA_17__7_, tempResultA_17__6_, tempResultA_17__5_, 
        tempResultA_17__4_, tempResultA_17__3_, tempResultA_17__2_, 
        tempResultA_17__1_, tempResultA_17__0_, tempResult[17]}), .cout(
        tempResultA_17__31_) );
  carryLookAheadAdder_14 generating_partialProducts_17__A1 ( .a({
        tempResultA_17__31_, tempResultA_17__30_, tempResultA_17__29_, 
        tempResultA_17__28_, tempResultA_17__27_, tempResultA_17__26_, 
        tempResultA_17__25_, tempResultA_17__24_, tempResultA_17__23_, 
        tempResultA_17__22_, tempResultA_17__21_, tempResultA_17__20_, 
        tempResultA_17__19_, tempResultA_17__18_, tempResultA_17__17_, 
        tempResultA_17__16_, tempResultA_17__15_, tempResultA_17__14_, 
        tempResultA_17__13_, tempResultA_17__12_, tempResultA_17__11_, 
        tempResultA_17__10_, tempResultA_17__9_, tempResultA_17__8_, 
        tempResultA_17__7_, tempResultA_17__6_, tempResultA_17__5_, 
        tempResultA_17__4_, tempResultA_17__3_, tempResultA_17__2_, 
        tempResultA_17__1_, tempResultA_17__0_}), .b(tempResultB[575:544]), 
        .cin(1'b0), .result({tempResultA_18__30_, tempResultA_18__29_, 
        tempResultA_18__28_, tempResultA_18__27_, tempResultA_18__26_, 
        tempResultA_18__25_, tempResultA_18__24_, tempResultA_18__23_, 
        tempResultA_18__22_, tempResultA_18__21_, tempResultA_18__20_, 
        tempResultA_18__19_, tempResultA_18__18_, tempResultA_18__17_, 
        tempResultA_18__16_, tempResultA_18__15_, tempResultA_18__14_, 
        tempResultA_18__13_, tempResultA_18__12_, tempResultA_18__11_, 
        tempResultA_18__10_, tempResultA_18__9_, tempResultA_18__8_, 
        tempResultA_18__7_, tempResultA_18__6_, tempResultA_18__5_, 
        tempResultA_18__4_, tempResultA_18__3_, tempResultA_18__2_, 
        tempResultA_18__1_, tempResultA_18__0_, tempResult[18]}), .cout(
        tempResultA_18__31_) );
  carryLookAheadAdder_13 generating_partialProducts_18__A1 ( .a({
        tempResultA_18__31_, tempResultA_18__30_, tempResultA_18__29_, 
        tempResultA_18__28_, tempResultA_18__27_, tempResultA_18__26_, 
        tempResultA_18__25_, tempResultA_18__24_, tempResultA_18__23_, 
        tempResultA_18__22_, tempResultA_18__21_, tempResultA_18__20_, 
        tempResultA_18__19_, tempResultA_18__18_, tempResultA_18__17_, 
        tempResultA_18__16_, tempResultA_18__15_, tempResultA_18__14_, 
        tempResultA_18__13_, tempResultA_18__12_, tempResultA_18__11_, 
        tempResultA_18__10_, tempResultA_18__9_, tempResultA_18__8_, 
        tempResultA_18__7_, tempResultA_18__6_, tempResultA_18__5_, 
        tempResultA_18__4_, tempResultA_18__3_, tempResultA_18__2_, 
        tempResultA_18__1_, tempResultA_18__0_}), .b(tempResultB[607:576]), 
        .cin(1'b0), .result({tempResultA_19__30_, tempResultA_19__29_, 
        tempResultA_19__28_, tempResultA_19__27_, tempResultA_19__26_, 
        tempResultA_19__25_, tempResultA_19__24_, tempResultA_19__23_, 
        tempResultA_19__22_, tempResultA_19__21_, tempResultA_19__20_, 
        tempResultA_19__19_, tempResultA_19__18_, tempResultA_19__17_, 
        tempResultA_19__16_, tempResultA_19__15_, tempResultA_19__14_, 
        tempResultA_19__13_, tempResultA_19__12_, tempResultA_19__11_, 
        tempResultA_19__10_, tempResultA_19__9_, tempResultA_19__8_, 
        tempResultA_19__7_, tempResultA_19__6_, tempResultA_19__5_, 
        tempResultA_19__4_, tempResultA_19__3_, tempResultA_19__2_, 
        tempResultA_19__1_, tempResultA_19__0_, tempResult[19]}), .cout(
        tempResultA_19__31_) );
  carryLookAheadAdder_12 generating_partialProducts_19__A1 ( .a({
        tempResultA_19__31_, tempResultA_19__30_, tempResultA_19__29_, 
        tempResultA_19__28_, tempResultA_19__27_, tempResultA_19__26_, 
        tempResultA_19__25_, tempResultA_19__24_, tempResultA_19__23_, 
        tempResultA_19__22_, tempResultA_19__21_, tempResultA_19__20_, 
        tempResultA_19__19_, tempResultA_19__18_, tempResultA_19__17_, 
        tempResultA_19__16_, tempResultA_19__15_, tempResultA_19__14_, 
        tempResultA_19__13_, tempResultA_19__12_, tempResultA_19__11_, 
        tempResultA_19__10_, tempResultA_19__9_, tempResultA_19__8_, 
        tempResultA_19__7_, tempResultA_19__6_, tempResultA_19__5_, 
        tempResultA_19__4_, tempResultA_19__3_, tempResultA_19__2_, 
        tempResultA_19__1_, tempResultA_19__0_}), .b(tempResultB[639:608]), 
        .cin(1'b0), .result({tempResultA_20__30_, tempResultA_20__29_, 
        tempResultA_20__28_, tempResultA_20__27_, tempResultA_20__26_, 
        tempResultA_20__25_, tempResultA_20__24_, tempResultA_20__23_, 
        tempResultA_20__22_, tempResultA_20__21_, tempResultA_20__20_, 
        tempResultA_20__19_, tempResultA_20__18_, tempResultA_20__17_, 
        tempResultA_20__16_, tempResultA_20__15_, tempResultA_20__14_, 
        tempResultA_20__13_, tempResultA_20__12_, tempResultA_20__11_, 
        tempResultA_20__10_, tempResultA_20__9_, tempResultA_20__8_, 
        tempResultA_20__7_, tempResultA_20__6_, tempResultA_20__5_, 
        tempResultA_20__4_, tempResultA_20__3_, tempResultA_20__2_, 
        tempResultA_20__1_, tempResultA_20__0_, tempResult[20]}), .cout(
        tempResultA_20__31_) );
  carryLookAheadAdder_11 generating_partialProducts_20__A1 ( .a({
        tempResultA_20__31_, tempResultA_20__30_, tempResultA_20__29_, 
        tempResultA_20__28_, tempResultA_20__27_, tempResultA_20__26_, 
        tempResultA_20__25_, tempResultA_20__24_, tempResultA_20__23_, 
        tempResultA_20__22_, tempResultA_20__21_, tempResultA_20__20_, 
        tempResultA_20__19_, tempResultA_20__18_, tempResultA_20__17_, 
        tempResultA_20__16_, tempResultA_20__15_, tempResultA_20__14_, 
        tempResultA_20__13_, tempResultA_20__12_, tempResultA_20__11_, 
        tempResultA_20__10_, tempResultA_20__9_, tempResultA_20__8_, 
        tempResultA_20__7_, tempResultA_20__6_, tempResultA_20__5_, 
        tempResultA_20__4_, tempResultA_20__3_, tempResultA_20__2_, 
        tempResultA_20__1_, tempResultA_20__0_}), .b(tempResultB[671:640]), 
        .cin(1'b0), .result({tempResultA_21__30_, tempResultA_21__29_, 
        tempResultA_21__28_, tempResultA_21__27_, tempResultA_21__26_, 
        tempResultA_21__25_, tempResultA_21__24_, tempResultA_21__23_, 
        tempResultA_21__22_, tempResultA_21__21_, tempResultA_21__20_, 
        tempResultA_21__19_, tempResultA_21__18_, tempResultA_21__17_, 
        tempResultA_21__16_, tempResultA_21__15_, tempResultA_21__14_, 
        tempResultA_21__13_, tempResultA_21__12_, tempResultA_21__11_, 
        tempResultA_21__10_, tempResultA_21__9_, tempResultA_21__8_, 
        tempResultA_21__7_, tempResultA_21__6_, tempResultA_21__5_, 
        tempResultA_21__4_, tempResultA_21__3_, tempResultA_21__2_, 
        tempResultA_21__1_, tempResultA_21__0_, tempResult[21]}), .cout(
        tempResultA_21__31_) );
  carryLookAheadAdder_10 generating_partialProducts_21__A1 ( .a({
        tempResultA_21__31_, tempResultA_21__30_, tempResultA_21__29_, 
        tempResultA_21__28_, tempResultA_21__27_, tempResultA_21__26_, 
        tempResultA_21__25_, tempResultA_21__24_, tempResultA_21__23_, 
        tempResultA_21__22_, tempResultA_21__21_, tempResultA_21__20_, 
        tempResultA_21__19_, tempResultA_21__18_, tempResultA_21__17_, 
        tempResultA_21__16_, tempResultA_21__15_, tempResultA_21__14_, 
        tempResultA_21__13_, tempResultA_21__12_, tempResultA_21__11_, 
        tempResultA_21__10_, tempResultA_21__9_, tempResultA_21__8_, 
        tempResultA_21__7_, tempResultA_21__6_, tempResultA_21__5_, 
        tempResultA_21__4_, tempResultA_21__3_, tempResultA_21__2_, 
        tempResultA_21__1_, tempResultA_21__0_}), .b(tempResultB[703:672]), 
        .cin(1'b0), .result({tempResultA_22__30_, tempResultA_22__29_, 
        tempResultA_22__28_, tempResultA_22__27_, tempResultA_22__26_, 
        tempResultA_22__25_, tempResultA_22__24_, tempResultA_22__23_, 
        tempResultA_22__22_, tempResultA_22__21_, tempResultA_22__20_, 
        tempResultA_22__19_, tempResultA_22__18_, tempResultA_22__17_, 
        tempResultA_22__16_, tempResultA_22__15_, tempResultA_22__14_, 
        tempResultA_22__13_, tempResultA_22__12_, tempResultA_22__11_, 
        tempResultA_22__10_, tempResultA_22__9_, tempResultA_22__8_, 
        tempResultA_22__7_, tempResultA_22__6_, tempResultA_22__5_, 
        tempResultA_22__4_, tempResultA_22__3_, tempResultA_22__2_, 
        tempResultA_22__1_, tempResultA_22__0_, tempResult[22]}), .cout(
        tempResultA_22__31_) );
  carryLookAheadAdder_9 generating_partialProducts_22__A1 ( .a({
        tempResultA_22__31_, tempResultA_22__30_, tempResultA_22__29_, 
        tempResultA_22__28_, tempResultA_22__27_, tempResultA_22__26_, 
        tempResultA_22__25_, tempResultA_22__24_, tempResultA_22__23_, 
        tempResultA_22__22_, tempResultA_22__21_, tempResultA_22__20_, 
        tempResultA_22__19_, tempResultA_22__18_, tempResultA_22__17_, 
        tempResultA_22__16_, tempResultA_22__15_, tempResultA_22__14_, 
        tempResultA_22__13_, tempResultA_22__12_, tempResultA_22__11_, 
        tempResultA_22__10_, tempResultA_22__9_, tempResultA_22__8_, 
        tempResultA_22__7_, tempResultA_22__6_, tempResultA_22__5_, 
        tempResultA_22__4_, tempResultA_22__3_, tempResultA_22__2_, 
        tempResultA_22__1_, tempResultA_22__0_}), .b(tempResultB[735:704]), 
        .cin(1'b0), .result({tempResultA_23__30_, tempResultA_23__29_, 
        tempResultA_23__28_, tempResultA_23__27_, tempResultA_23__26_, 
        tempResultA_23__25_, tempResultA_23__24_, tempResultA_23__23_, 
        tempResultA_23__22_, tempResultA_23__21_, tempResultA_23__20_, 
        tempResultA_23__19_, tempResultA_23__18_, tempResultA_23__17_, 
        tempResultA_23__16_, tempResultA_23__15_, tempResultA_23__14_, 
        tempResultA_23__13_, tempResultA_23__12_, tempResultA_23__11_, 
        tempResultA_23__10_, tempResultA_23__9_, tempResultA_23__8_, 
        tempResultA_23__7_, tempResultA_23__6_, tempResultA_23__5_, 
        tempResultA_23__4_, tempResultA_23__3_, tempResultA_23__2_, 
        tempResultA_23__1_, tempResultA_23__0_, tempResult[23]}), .cout(
        tempResultA_23__31_) );
  carryLookAheadAdder_8 generating_partialProducts_23__A1 ( .a({
        tempResultA_23__31_, tempResultA_23__30_, tempResultA_23__29_, 
        tempResultA_23__28_, tempResultA_23__27_, tempResultA_23__26_, 
        tempResultA_23__25_, tempResultA_23__24_, tempResultA_23__23_, 
        tempResultA_23__22_, tempResultA_23__21_, tempResultA_23__20_, 
        tempResultA_23__19_, tempResultA_23__18_, tempResultA_23__17_, 
        tempResultA_23__16_, tempResultA_23__15_, tempResultA_23__14_, 
        tempResultA_23__13_, tempResultA_23__12_, tempResultA_23__11_, 
        tempResultA_23__10_, tempResultA_23__9_, tempResultA_23__8_, 
        tempResultA_23__7_, tempResultA_23__6_, tempResultA_23__5_, 
        tempResultA_23__4_, tempResultA_23__3_, tempResultA_23__2_, 
        tempResultA_23__1_, tempResultA_23__0_}), .b(tempResultB[767:736]), 
        .cin(1'b0), .result({tempResultA_24__30_, tempResultA_24__29_, 
        tempResultA_24__28_, tempResultA_24__27_, tempResultA_24__26_, 
        tempResultA_24__25_, tempResultA_24__24_, tempResultA_24__23_, 
        tempResultA_24__22_, tempResultA_24__21_, tempResultA_24__20_, 
        tempResultA_24__19_, tempResultA_24__18_, tempResultA_24__17_, 
        tempResultA_24__16_, tempResultA_24__15_, tempResultA_24__14_, 
        tempResultA_24__13_, tempResultA_24__12_, tempResultA_24__11_, 
        tempResultA_24__10_, tempResultA_24__9_, tempResultA_24__8_, 
        tempResultA_24__7_, tempResultA_24__6_, tempResultA_24__5_, 
        tempResultA_24__4_, tempResultA_24__3_, tempResultA_24__2_, 
        tempResultA_24__1_, tempResultA_24__0_, tempResult[24]}), .cout(
        tempResultA_24__31_) );
  carryLookAheadAdder_7 generating_partialProducts_24__A1 ( .a({
        tempResultA_24__31_, tempResultA_24__30_, tempResultA_24__29_, 
        tempResultA_24__28_, tempResultA_24__27_, tempResultA_24__26_, 
        tempResultA_24__25_, tempResultA_24__24_, tempResultA_24__23_, 
        tempResultA_24__22_, tempResultA_24__21_, tempResultA_24__20_, 
        tempResultA_24__19_, tempResultA_24__18_, tempResultA_24__17_, 
        tempResultA_24__16_, tempResultA_24__15_, tempResultA_24__14_, 
        tempResultA_24__13_, tempResultA_24__12_, tempResultA_24__11_, 
        tempResultA_24__10_, tempResultA_24__9_, tempResultA_24__8_, 
        tempResultA_24__7_, tempResultA_24__6_, tempResultA_24__5_, 
        tempResultA_24__4_, tempResultA_24__3_, tempResultA_24__2_, 
        tempResultA_24__1_, tempResultA_24__0_}), .b(tempResultB[799:768]), 
        .cin(1'b0), .result({tempResultA_25__30_, tempResultA_25__29_, 
        tempResultA_25__28_, tempResultA_25__27_, tempResultA_25__26_, 
        tempResultA_25__25_, tempResultA_25__24_, tempResultA_25__23_, 
        tempResultA_25__22_, tempResultA_25__21_, tempResultA_25__20_, 
        tempResultA_25__19_, tempResultA_25__18_, tempResultA_25__17_, 
        tempResultA_25__16_, tempResultA_25__15_, tempResultA_25__14_, 
        tempResultA_25__13_, tempResultA_25__12_, tempResultA_25__11_, 
        tempResultA_25__10_, tempResultA_25__9_, tempResultA_25__8_, 
        tempResultA_25__7_, tempResultA_25__6_, tempResultA_25__5_, 
        tempResultA_25__4_, tempResultA_25__3_, tempResultA_25__2_, 
        tempResultA_25__1_, tempResultA_25__0_, tempResult[25]}), .cout(
        tempResultA_25__31_) );
  carryLookAheadAdder_6 generating_partialProducts_25__A1 ( .a({
        tempResultA_25__31_, tempResultA_25__30_, tempResultA_25__29_, 
        tempResultA_25__28_, tempResultA_25__27_, tempResultA_25__26_, 
        tempResultA_25__25_, tempResultA_25__24_, tempResultA_25__23_, 
        tempResultA_25__22_, tempResultA_25__21_, tempResultA_25__20_, 
        tempResultA_25__19_, tempResultA_25__18_, tempResultA_25__17_, 
        tempResultA_25__16_, tempResultA_25__15_, tempResultA_25__14_, 
        tempResultA_25__13_, tempResultA_25__12_, tempResultA_25__11_, 
        tempResultA_25__10_, tempResultA_25__9_, tempResultA_25__8_, 
        tempResultA_25__7_, tempResultA_25__6_, tempResultA_25__5_, 
        tempResultA_25__4_, tempResultA_25__3_, tempResultA_25__2_, 
        tempResultA_25__1_, tempResultA_25__0_}), .b(tempResultB[831:800]), 
        .cin(1'b0), .result({tempResultA_26__30_, tempResultA_26__29_, 
        tempResultA_26__28_, tempResultA_26__27_, tempResultA_26__26_, 
        tempResultA_26__25_, tempResultA_26__24_, tempResultA_26__23_, 
        tempResultA_26__22_, tempResultA_26__21_, tempResultA_26__20_, 
        tempResultA_26__19_, tempResultA_26__18_, tempResultA_26__17_, 
        tempResultA_26__16_, tempResultA_26__15_, tempResultA_26__14_, 
        tempResultA_26__13_, tempResultA_26__12_, tempResultA_26__11_, 
        tempResultA_26__10_, tempResultA_26__9_, tempResultA_26__8_, 
        tempResultA_26__7_, tempResultA_26__6_, tempResultA_26__5_, 
        tempResultA_26__4_, tempResultA_26__3_, tempResultA_26__2_, 
        tempResultA_26__1_, tempResultA_26__0_, tempResult[26]}), .cout(
        tempResultA_26__31_) );
  carryLookAheadAdder_5 generating_partialProducts_26__A1 ( .a({
        tempResultA_26__31_, tempResultA_26__30_, tempResultA_26__29_, 
        tempResultA_26__28_, tempResultA_26__27_, tempResultA_26__26_, 
        tempResultA_26__25_, tempResultA_26__24_, tempResultA_26__23_, 
        tempResultA_26__22_, tempResultA_26__21_, tempResultA_26__20_, 
        tempResultA_26__19_, tempResultA_26__18_, tempResultA_26__17_, 
        tempResultA_26__16_, tempResultA_26__15_, tempResultA_26__14_, 
        tempResultA_26__13_, tempResultA_26__12_, tempResultA_26__11_, 
        tempResultA_26__10_, tempResultA_26__9_, tempResultA_26__8_, 
        tempResultA_26__7_, tempResultA_26__6_, tempResultA_26__5_, 
        tempResultA_26__4_, tempResultA_26__3_, tempResultA_26__2_, 
        tempResultA_26__1_, tempResultA_26__0_}), .b(tempResultB[863:832]), 
        .cin(1'b0), .result({tempResultA_27__30_, tempResultA_27__29_, 
        tempResultA_27__28_, tempResultA_27__27_, tempResultA_27__26_, 
        tempResultA_27__25_, tempResultA_27__24_, tempResultA_27__23_, 
        tempResultA_27__22_, tempResultA_27__21_, tempResultA_27__20_, 
        tempResultA_27__19_, tempResultA_27__18_, tempResultA_27__17_, 
        tempResultA_27__16_, tempResultA_27__15_, tempResultA_27__14_, 
        tempResultA_27__13_, tempResultA_27__12_, tempResultA_27__11_, 
        tempResultA_27__10_, tempResultA_27__9_, tempResultA_27__8_, 
        tempResultA_27__7_, tempResultA_27__6_, tempResultA_27__5_, 
        tempResultA_27__4_, tempResultA_27__3_, tempResultA_27__2_, 
        tempResultA_27__1_, tempResultA_27__0_, tempResult[27]}), .cout(
        tempResultA_27__31_) );
  carryLookAheadAdder_4 generating_partialProducts_27__A1 ( .a({
        tempResultA_27__31_, tempResultA_27__30_, tempResultA_27__29_, 
        tempResultA_27__28_, tempResultA_27__27_, tempResultA_27__26_, 
        tempResultA_27__25_, tempResultA_27__24_, tempResultA_27__23_, 
        tempResultA_27__22_, tempResultA_27__21_, tempResultA_27__20_, 
        tempResultA_27__19_, tempResultA_27__18_, tempResultA_27__17_, 
        tempResultA_27__16_, tempResultA_27__15_, tempResultA_27__14_, 
        tempResultA_27__13_, tempResultA_27__12_, tempResultA_27__11_, 
        tempResultA_27__10_, tempResultA_27__9_, tempResultA_27__8_, 
        tempResultA_27__7_, tempResultA_27__6_, tempResultA_27__5_, 
        tempResultA_27__4_, tempResultA_27__3_, tempResultA_27__2_, 
        tempResultA_27__1_, tempResultA_27__0_}), .b(tempResultB[895:864]), 
        .cin(1'b0), .result({tempResultA_28__30_, tempResultA_28__29_, 
        tempResultA_28__28_, tempResultA_28__27_, tempResultA_28__26_, 
        tempResultA_28__25_, tempResultA_28__24_, tempResultA_28__23_, 
        tempResultA_28__22_, tempResultA_28__21_, tempResultA_28__20_, 
        tempResultA_28__19_, tempResultA_28__18_, tempResultA_28__17_, 
        tempResultA_28__16_, tempResultA_28__15_, tempResultA_28__14_, 
        tempResultA_28__13_, tempResultA_28__12_, tempResultA_28__11_, 
        tempResultA_28__10_, tempResultA_28__9_, tempResultA_28__8_, 
        tempResultA_28__7_, tempResultA_28__6_, tempResultA_28__5_, 
        tempResultA_28__4_, tempResultA_28__3_, tempResultA_28__2_, 
        tempResultA_28__1_, tempResultA_28__0_, tempResult[28]}), .cout(
        tempResultA_28__31_) );
  carryLookAheadAdder_3 generating_partialProducts_28__A1 ( .a({
        tempResultA_28__31_, tempResultA_28__30_, tempResultA_28__29_, 
        tempResultA_28__28_, tempResultA_28__27_, tempResultA_28__26_, 
        tempResultA_28__25_, tempResultA_28__24_, tempResultA_28__23_, 
        tempResultA_28__22_, tempResultA_28__21_, tempResultA_28__20_, 
        tempResultA_28__19_, tempResultA_28__18_, tempResultA_28__17_, 
        tempResultA_28__16_, tempResultA_28__15_, tempResultA_28__14_, 
        tempResultA_28__13_, tempResultA_28__12_, tempResultA_28__11_, 
        tempResultA_28__10_, tempResultA_28__9_, tempResultA_28__8_, 
        tempResultA_28__7_, tempResultA_28__6_, tempResultA_28__5_, 
        tempResultA_28__4_, tempResultA_28__3_, tempResultA_28__2_, 
        tempResultA_28__1_, tempResultA_28__0_}), .b(tempResultB[927:896]), 
        .cin(1'b0), .result({tempResultA_29__30_, tempResultA_29__29_, 
        tempResultA_29__28_, tempResultA_29__27_, tempResultA_29__26_, 
        tempResultA_29__25_, tempResultA_29__24_, tempResultA_29__23_, 
        tempResultA_29__22_, tempResultA_29__21_, tempResultA_29__20_, 
        tempResultA_29__19_, tempResultA_29__18_, tempResultA_29__17_, 
        tempResultA_29__16_, tempResultA_29__15_, tempResultA_29__14_, 
        tempResultA_29__13_, tempResultA_29__12_, tempResultA_29__11_, 
        tempResultA_29__10_, tempResultA_29__9_, tempResultA_29__8_, 
        tempResultA_29__7_, tempResultA_29__6_, tempResultA_29__5_, 
        tempResultA_29__4_, tempResultA_29__3_, tempResultA_29__2_, 
        tempResultA_29__1_, tempResultA_29__0_, tempResult[29]}), .cout(
        tempResultA_29__31_) );
  carryLookAheadAdder_2 generating_partialProducts_29__A1 ( .a({
        tempResultA_29__31_, tempResultA_29__30_, tempResultA_29__29_, 
        tempResultA_29__28_, tempResultA_29__27_, tempResultA_29__26_, 
        tempResultA_29__25_, tempResultA_29__24_, tempResultA_29__23_, 
        tempResultA_29__22_, tempResultA_29__21_, tempResultA_29__20_, 
        tempResultA_29__19_, tempResultA_29__18_, tempResultA_29__17_, 
        tempResultA_29__16_, tempResultA_29__15_, tempResultA_29__14_, 
        tempResultA_29__13_, tempResultA_29__12_, tempResultA_29__11_, 
        tempResultA_29__10_, tempResultA_29__9_, tempResultA_29__8_, 
        tempResultA_29__7_, tempResultA_29__6_, tempResultA_29__5_, 
        tempResultA_29__4_, tempResultA_29__3_, tempResultA_29__2_, 
        tempResultA_29__1_, tempResultA_29__0_}), .b(tempResultB[959:928]), 
        .cin(1'b0), .result({tempResultA_30__30_, tempResultA_30__29_, 
        tempResultA_30__28_, tempResultA_30__27_, tempResultA_30__26_, 
        tempResultA_30__25_, tempResultA_30__24_, tempResultA_30__23_, 
        tempResultA_30__22_, tempResultA_30__21_, tempResultA_30__20_, 
        tempResultA_30__19_, tempResultA_30__18_, tempResultA_30__17_, 
        tempResultA_30__16_, tempResultA_30__15_, tempResultA_30__14_, 
        tempResultA_30__13_, tempResultA_30__12_, tempResultA_30__11_, 
        tempResultA_30__10_, tempResultA_30__9_, tempResultA_30__8_, 
        tempResultA_30__7_, tempResultA_30__6_, tempResultA_30__5_, 
        tempResultA_30__4_, tempResultA_30__3_, tempResultA_30__2_, 
        tempResultA_30__1_, tempResultA_30__0_, tempResult[30]}), .cout(
        tempResultA_30__31_) );
  carryLookAheadAdder_1 A2 ( .a({tempResultA_30__31_, tempResultA_30__30_, 
        tempResultA_30__29_, tempResultA_30__28_, tempResultA_30__27_, 
        tempResultA_30__26_, tempResultA_30__25_, tempResultA_30__24_, 
        tempResultA_30__23_, tempResultA_30__22_, tempResultA_30__21_, 
        tempResultA_30__20_, tempResultA_30__19_, tempResultA_30__18_, 
        tempResultA_30__17_, tempResultA_30__16_, tempResultA_30__15_, 
        tempResultA_30__14_, tempResultA_30__13_, tempResultA_30__12_, 
        tempResultA_30__11_, tempResultA_30__10_, tempResultA_30__9_, 
        tempResultA_30__8_, tempResultA_30__7_, tempResultA_30__6_, 
        tempResultA_30__5_, tempResultA_30__4_, tempResultA_30__3_, 
        tempResultA_30__2_, tempResultA_30__1_, tempResultA_30__0_}), .b(
        tempResultB[991:960]), .cin(1'b0), .result(tempResult[62:31]), .cout(
        tempResult[63]) );
  multiplierTreeV2_DW01_add_0 add_32 ( .A({N62, N63, N64, N65, N66, N67, N68, 
        N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, 
        N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, 
        N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, 
        N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, 
        N121, N122, N123, N124, N125}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n193}), .CI(1'b0), .SUM(result) );
  multiplierTreeV2_DW01_add_1 add_15 ( .A({1'b0, N31, N32, N33, N34, N35, N36, 
        N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, 
        N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n197}), .CI(1'b0), .SUM(b_abs) );
  multiplierTreeV2_DW01_add_2 add_14 ( .A({1'b0, N0, N1, N2, N3, N4, N5, N6, 
        N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, 
        N22, N23, N24, N25, N26, N27, N28, N29, N30}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, n199}), .CI(1'b0), .SUM(a_abs) );
  BUF_X1 U5 ( .A(n260), .Z(n180) );
  NOR2_X1 U6 ( .A1(n38), .A2(n161), .ZN(tempResultB[274]) );
  NOR2_X1 U7 ( .A1(n28), .A2(n168), .ZN(tempResultB[214]) );
  NOR2_X1 U8 ( .A1(n32), .A2(n162), .ZN(tempResultB[276]) );
  NOR2_X1 U9 ( .A1(n26), .A2(n168), .ZN(tempResultB[215]) );
  NOR2_X1 U10 ( .A1(n20), .A2(n174), .ZN(tempResultB[154]) );
  NOR2_X1 U11 ( .A1(n28), .A2(n162), .ZN(tempResultB[278]) );
  NOR2_X1 U12 ( .A1(n59), .A2(n137), .ZN(tempResultB[523]) );
  NOR2_X1 U13 ( .A1(n59), .A2(n134), .ZN(tempResultB[555]) );
  NOR2_X1 U14 ( .A1(n59), .A2(n131), .ZN(tempResultB[587]) );
  NOR2_X1 U15 ( .A1(n65), .A2(n133), .ZN(tempResultB[585]) );
  NOR2_X1 U16 ( .A1(n65), .A2(n127), .ZN(tempResultB[649]) );
  NOR2_X1 U17 ( .A1(n72), .A2(n115), .ZN(tempResultB[775]) );
  NOR2_X1 U18 ( .A1(n78), .A2(n130), .ZN(tempResultB[613]) );
  BUF_X1 U19 ( .A(n220), .Z(n59) );
  BUF_X1 U20 ( .A(n227), .Z(n82) );
  NOR2_X1 U21 ( .A1(n83), .A2(n103), .ZN(tempResultB[899]) );
  NOR2_X1 U22 ( .A1(n67), .A2(n103), .ZN(tempResultB[904]) );
  BUF_X1 U23 ( .A(n201), .Z(n13) );
  INV_X1 U24 ( .A(b_abs[2]), .ZN(n261) );
  INV_X1 U25 ( .A(b_abs[3]), .ZN(n260) );
  INV_X1 U26 ( .A(b_abs[4]), .ZN(n259) );
  INV_X1 U27 ( .A(b_abs[5]), .ZN(n258) );
  INV_X1 U28 ( .A(b_abs[6]), .ZN(n257) );
  INV_X1 U29 ( .A(b_abs[7]), .ZN(n256) );
  INV_X1 U30 ( .A(b_abs[8]), .ZN(n255) );
  INV_X1 U31 ( .A(b_abs[9]), .ZN(n254) );
  INV_X1 U32 ( .A(b_abs[10]), .ZN(n253) );
  INV_X1 U33 ( .A(b_abs[11]), .ZN(n252) );
  INV_X1 U34 ( .A(b_abs[12]), .ZN(n251) );
  INV_X1 U35 ( .A(b_abs[13]), .ZN(n250) );
  INV_X1 U36 ( .A(b_abs[14]), .ZN(n249) );
  INV_X1 U37 ( .A(b_abs[15]), .ZN(n248) );
  INV_X1 U38 ( .A(b_abs[16]), .ZN(n247) );
  INV_X1 U39 ( .A(b_abs[17]), .ZN(n246) );
  INV_X1 U40 ( .A(b_abs[18]), .ZN(n245) );
  INV_X1 U41 ( .A(b_abs[19]), .ZN(n244) );
  INV_X1 U42 ( .A(b_abs[20]), .ZN(n243) );
  INV_X1 U43 ( .A(b_abs[21]), .ZN(n242) );
  INV_X1 U44 ( .A(b_abs[22]), .ZN(n241) );
  INV_X1 U45 ( .A(b_abs[23]), .ZN(n240) );
  INV_X1 U46 ( .A(b_abs[24]), .ZN(n239) );
  INV_X1 U47 ( .A(b_abs[25]), .ZN(n238) );
  INV_X1 U48 ( .A(b_abs[26]), .ZN(n237) );
  INV_X1 U49 ( .A(b_abs[27]), .ZN(n236) );
  INV_X1 U50 ( .A(b_abs[28]), .ZN(n235) );
  INV_X1 U51 ( .A(a_abs[1]), .ZN(n230) );
  INV_X1 U52 ( .A(a_abs[2]), .ZN(n229) );
  INV_X1 U53 ( .A(a_abs[3]), .ZN(n228) );
  NOR2_X1 U54 ( .A1(n77), .A2(n100), .ZN(tempResultB[933]) );
  INV_X1 U55 ( .A(a_abs[5]), .ZN(n226) );
  INV_X1 U56 ( .A(a_abs[6]), .ZN(n225) );
  INV_X1 U57 ( .A(a_abs[8]), .ZN(n223) );
  INV_X1 U58 ( .A(a_abs[10]), .ZN(n221) );
  INV_X1 U59 ( .A(a_abs[12]), .ZN(n219) );
  INV_X1 U60 ( .A(a_abs[13]), .ZN(n218) );
  INV_X1 U61 ( .A(a_abs[15]), .ZN(n216) );
  INV_X1 U62 ( .A(a_abs[16]), .ZN(n215) );
  INV_X1 U63 ( .A(a_abs[17]), .ZN(n214) );
  INV_X1 U64 ( .A(a_abs[28]), .ZN(n203) );
  INV_X1 U65 ( .A(b_abs[29]), .ZN(n234) );
  BUF_X1 U66 ( .A(n261), .Z(n182) );
  INV_X1 U67 ( .A(b_abs[30]), .ZN(n233) );
  INV_X1 U68 ( .A(a_abs[31]), .ZN(n200) );
  INV_X1 U69 ( .A(b_abs[31]), .ZN(n232) );
  BUF_X1 U70 ( .A(n201), .Z(n12) );
  INV_X1 U71 ( .A(a_abs[0]), .ZN(n231) );
  BUF_X1 U72 ( .A(n191), .Z(n193) );
  CLKBUF_X1 U73 ( .A(n262), .Z(n187) );
  BUF_X1 U74 ( .A(n222), .Z(n65) );
  BUF_X1 U75 ( .A(n213), .Z(n39) );
  BUF_X1 U76 ( .A(n208), .Z(n27) );
  BUF_X1 U77 ( .A(n224), .Z(n72) );
  BUF_X1 U78 ( .A(n226), .Z(n78) );
  BUF_X1 U79 ( .A(n211), .Z(n33) );
  BUF_X1 U80 ( .A(n214), .Z(n41) );
  BUF_X1 U81 ( .A(n215), .Z(n44) );
  BUF_X1 U82 ( .A(n219), .Z(n56) );
  BUF_X1 U83 ( .A(n218), .Z(n53) );
  BUF_X1 U84 ( .A(n216), .Z(n47) );
  BUF_X1 U85 ( .A(n217), .Z(n50) );
  BUF_X1 U86 ( .A(n212), .Z(n36) );
  BUF_X1 U87 ( .A(n221), .Z(n62) );
  BUF_X1 U88 ( .A(n228), .Z(n84) );
  BUF_X1 U89 ( .A(n227), .Z(n81) );
  BUF_X1 U90 ( .A(n223), .Z(n69) );
  BUF_X1 U91 ( .A(n225), .Z(n75) );
  BUF_X1 U92 ( .A(n230), .Z(n90) );
  BUF_X1 U93 ( .A(n229), .Z(n87) );
  BUF_X1 U94 ( .A(n231), .Z(n93) );
  BUF_X1 U95 ( .A(n261), .Z(n183) );
  BUF_X1 U96 ( .A(n259), .Z(n176) );
  BUF_X1 U97 ( .A(n260), .Z(n179) );
  BUF_X1 U98 ( .A(n200), .Z(n11) );
  BUF_X1 U99 ( .A(n218), .Z(n54) );
  BUF_X1 U100 ( .A(n261), .Z(n184) );
  BUF_X1 U101 ( .A(n260), .Z(n181) );
  BUF_X1 U102 ( .A(n209), .Z(n28) );
  BUF_X1 U103 ( .A(n205), .Z(n20) );
  BUF_X1 U104 ( .A(n202), .Z(n14) );
  BUF_X1 U105 ( .A(n203), .Z(n16) );
  BUF_X1 U106 ( .A(n204), .Z(n18) );
  BUF_X1 U107 ( .A(n207), .Z(n24) );
  BUF_X1 U108 ( .A(n206), .Z(n22) );
  BUF_X1 U109 ( .A(n200), .Z(n10) );
  XOR2_X1 U110 ( .A(n8), .B(a[1]), .Z(N29) );
  CLKBUF_X1 U111 ( .A(n262), .Z(n185) );
  NOR2_X1 U112 ( .A1(n38), .A2(n179), .ZN(tempResultB[82]) );
  NOR2_X1 U113 ( .A1(n26), .A2(n180), .ZN(tempResultB[87]) );
  NOR2_X1 U114 ( .A1(n38), .A2(n176), .ZN(tempResultB[114]) );
  NOR2_X1 U115 ( .A1(n38), .A2(n173), .ZN(tempResultB[146]) );
  NOR2_X1 U116 ( .A1(n38), .A2(n170), .ZN(tempResultB[178]) );
  NOR2_X1 U117 ( .A1(n26), .A2(n177), .ZN(tempResultB[119]) );
  NOR2_X1 U118 ( .A1(n38), .A2(n167), .ZN(tempResultB[210]) );
  NOR2_X1 U119 ( .A1(n26), .A2(n174), .ZN(tempResultB[151]) );
  NOR2_X1 U120 ( .A1(n26), .A2(n171), .ZN(tempResultB[183]) );
  XOR2_X1 U121 ( .A(tempResult[34]), .B(n193), .Z(N91) );
  NOR2_X1 U122 ( .A1(n32), .A2(n180), .ZN(tempResultB[84]) );
  NOR2_X1 U123 ( .A1(n32), .A2(n177), .ZN(tempResultB[116]) );
  NOR2_X1 U124 ( .A1(n32), .A2(n174), .ZN(tempResultB[148]) );
  NOR2_X1 U125 ( .A1(n32), .A2(n171), .ZN(tempResultB[180]) );
  NOR2_X1 U126 ( .A1(n31), .A2(n183), .ZN(tempResultB[53]) );
  NOR2_X1 U127 ( .A1(n15), .A2(n183), .ZN(tempResultB[61]) );
  NOR2_X1 U128 ( .A1(n29), .A2(n183), .ZN(tempResultB[54]) );
  NOR2_X1 U129 ( .A1(n19), .A2(n183), .ZN(tempResultB[59]) );
  NOR2_X1 U130 ( .A1(n23), .A2(n183), .ZN(tempResultB[57]) );
  NOR2_X1 U131 ( .A1(n11), .A2(n190), .ZN(tempResultA_0__30_) );
  NOR2_X1 U132 ( .A1(n91), .A2(n188), .ZN(tempResultA_0__0_) );
  NOR2_X1 U133 ( .A1(n11), .A2(n187), .ZN(tempResultB[31]) );
  NOR2_X1 U134 ( .A1(n13), .A2(n183), .ZN(tempResultB[62]) );
  NOR2_X1 U135 ( .A1(n94), .A2(n262), .ZN(tempResultB[0]) );
  NOR2_X1 U136 ( .A1(n12), .A2(n180), .ZN(tempResultB[94]) );
  NOR2_X1 U137 ( .A1(n12), .A2(n177), .ZN(tempResultB[126]) );
  NOR2_X1 U138 ( .A1(n12), .A2(n174), .ZN(tempResultB[158]) );
  NOR2_X1 U139 ( .A1(n12), .A2(n171), .ZN(tempResultB[190]) );
  NOR2_X1 U140 ( .A1(n10), .A2(n184), .ZN(tempResultB[63]) );
  NOR2_X1 U141 ( .A1(n9), .A2(n181), .ZN(tempResultB[95]) );
  NOR2_X1 U142 ( .A1(n9), .A2(n178), .ZN(tempResultB[127]) );
  NOR2_X1 U143 ( .A1(n9), .A2(n175), .ZN(tempResultB[159]) );
  NOR2_X1 U144 ( .A1(n9), .A2(n172), .ZN(tempResultB[191]) );
  NOR2_X1 U145 ( .A1(n93), .A2(n182), .ZN(tempResultB[32]) );
  NOR2_X1 U146 ( .A1(n92), .A2(n176), .ZN(tempResultB[96]) );
  NOR2_X1 U147 ( .A1(n92), .A2(n179), .ZN(tempResultB[64]) );
  NOR2_X1 U148 ( .A1(n92), .A2(n173), .ZN(tempResultB[128]) );
  NOR2_X1 U149 ( .A1(n92), .A2(n170), .ZN(tempResultB[160]) );
  NOR2_X1 U150 ( .A1(n92), .A2(n167), .ZN(tempResultB[192]) );
  NOR2_X1 U151 ( .A1(n92), .A2(n164), .ZN(tempResultB[224]) );
  NOR2_X1 U152 ( .A1(n92), .A2(n161), .ZN(tempResultB[256]) );
  NOR2_X1 U153 ( .A1(n58), .A2(n179), .ZN(tempResultB[75]) );
  NOR2_X1 U154 ( .A1(n58), .A2(n176), .ZN(tempResultB[107]) );
  NOR2_X1 U155 ( .A1(n58), .A2(n173), .ZN(tempResultB[139]) );
  NOR2_X1 U156 ( .A1(n58), .A2(n170), .ZN(tempResultB[171]) );
  NOR2_X1 U157 ( .A1(n59), .A2(n182), .ZN(tempResultB[43]) );
  NOR2_X1 U158 ( .A1(n25), .A2(n183), .ZN(tempResultB[56]) );
  NOR2_X1 U159 ( .A1(n91), .A2(n262), .ZN(tempResultB[1]) );
  NOR2_X1 U160 ( .A1(n83), .A2(n181), .ZN(tempResultB[67]) );
  NOR2_X1 U161 ( .A1(n84), .A2(n184), .ZN(tempResultB[35]) );
  NOR2_X1 U162 ( .A1(n65), .A2(n184), .ZN(tempResultB[41]) );
  NOR2_X1 U163 ( .A1(n81), .A2(n184), .ZN(tempResultB[36]) );
  NOR2_X1 U164 ( .A1(n69), .A2(n184), .ZN(tempResultB[40]) );
  NOR2_X1 U165 ( .A1(n72), .A2(n184), .ZN(tempResultB[39]) );
  NOR2_X1 U166 ( .A1(n75), .A2(n184), .ZN(tempResultB[38]) );
  NOR2_X1 U167 ( .A1(n78), .A2(n184), .ZN(tempResultB[37]) );
  NOR2_X1 U168 ( .A1(n80), .A2(n181), .ZN(tempResultB[68]) );
  NOR2_X1 U169 ( .A1(n77), .A2(n181), .ZN(tempResultB[69]) );
  NOR2_X1 U170 ( .A1(n83), .A2(n178), .ZN(tempResultB[99]) );
  NOR2_X1 U171 ( .A1(n74), .A2(n181), .ZN(tempResultB[70]) );
  NOR2_X1 U172 ( .A1(n80), .A2(n178), .ZN(tempResultB[100]) );
  NOR2_X1 U173 ( .A1(n71), .A2(n181), .ZN(tempResultB[71]) );
  NOR2_X1 U174 ( .A1(n77), .A2(n178), .ZN(tempResultB[101]) );
  NOR2_X1 U175 ( .A1(n83), .A2(n175), .ZN(tempResultB[131]) );
  NOR2_X1 U176 ( .A1(n67), .A2(n181), .ZN(tempResultB[72]) );
  NOR2_X1 U177 ( .A1(n74), .A2(n178), .ZN(tempResultB[102]) );
  NOR2_X1 U178 ( .A1(n80), .A2(n175), .ZN(tempResultB[132]) );
  NOR2_X1 U179 ( .A1(n71), .A2(n178), .ZN(tempResultB[103]) );
  NOR2_X1 U180 ( .A1(n77), .A2(n175), .ZN(tempResultB[133]) );
  NOR2_X1 U181 ( .A1(n83), .A2(n172), .ZN(tempResultB[163]) );
  NOR2_X1 U182 ( .A1(n64), .A2(n181), .ZN(tempResultB[73]) );
  NOR2_X1 U183 ( .A1(n67), .A2(n178), .ZN(tempResultB[104]) );
  NOR2_X1 U184 ( .A1(n74), .A2(n175), .ZN(tempResultB[134]) );
  NOR2_X1 U185 ( .A1(n80), .A2(n172), .ZN(tempResultB[164]) );
  NOR2_X1 U186 ( .A1(n71), .A2(n175), .ZN(tempResultB[135]) );
  NOR2_X1 U187 ( .A1(n77), .A2(n172), .ZN(tempResultB[165]) );
  NOR2_X1 U188 ( .A1(n83), .A2(n169), .ZN(tempResultB[195]) );
  NOR2_X1 U189 ( .A1(n64), .A2(n178), .ZN(tempResultB[105]) );
  NOR2_X1 U190 ( .A1(n67), .A2(n175), .ZN(tempResultB[136]) );
  NOR2_X1 U191 ( .A1(n74), .A2(n172), .ZN(tempResultB[166]) );
  NOR2_X1 U192 ( .A1(n80), .A2(n169), .ZN(tempResultB[196]) );
  NOR2_X1 U193 ( .A1(n71), .A2(n172), .ZN(tempResultB[167]) );
  NOR2_X1 U194 ( .A1(n77), .A2(n169), .ZN(tempResultB[197]) );
  NOR2_X1 U195 ( .A1(n83), .A2(n166), .ZN(tempResultB[227]) );
  NOR2_X1 U196 ( .A1(n64), .A2(n175), .ZN(tempResultB[137]) );
  NOR2_X1 U197 ( .A1(n67), .A2(n172), .ZN(tempResultB[168]) );
  NOR2_X1 U198 ( .A1(n64), .A2(n172), .ZN(tempResultB[169]) );
  NOR2_X1 U199 ( .A1(n14), .A2(n180), .ZN(tempResultB[93]) );
  NOR2_X1 U200 ( .A1(n16), .A2(n180), .ZN(tempResultB[92]) );
  NOR2_X1 U201 ( .A1(n28), .A2(n180), .ZN(tempResultB[86]) );
  NOR2_X1 U202 ( .A1(n18), .A2(n180), .ZN(tempResultB[91]) );
  NOR2_X1 U203 ( .A1(n20), .A2(n180), .ZN(tempResultB[90]) );
  NOR2_X1 U204 ( .A1(n24), .A2(n180), .ZN(tempResultB[88]) );
  NOR2_X1 U205 ( .A1(n22), .A2(n180), .ZN(tempResultB[89]) );
  NOR2_X1 U206 ( .A1(n30), .A2(n180), .ZN(tempResultB[85]) );
  NOR2_X1 U207 ( .A1(n30), .A2(n177), .ZN(tempResultB[117]) );
  NOR2_X1 U208 ( .A1(n28), .A2(n177), .ZN(tempResultB[118]) );
  NOR2_X1 U209 ( .A1(n30), .A2(n174), .ZN(tempResultB[149]) );
  NOR2_X1 U210 ( .A1(n24), .A2(n177), .ZN(tempResultB[120]) );
  NOR2_X1 U211 ( .A1(n28), .A2(n174), .ZN(tempResultB[150]) );
  NOR2_X1 U212 ( .A1(n22), .A2(n177), .ZN(tempResultB[121]) );
  NOR2_X1 U213 ( .A1(n30), .A2(n171), .ZN(tempResultB[181]) );
  NOR2_X1 U214 ( .A1(n20), .A2(n177), .ZN(tempResultB[122]) );
  NOR2_X1 U215 ( .A1(n24), .A2(n174), .ZN(tempResultB[152]) );
  NOR2_X1 U216 ( .A1(n28), .A2(n171), .ZN(tempResultB[182]) );
  NOR2_X1 U217 ( .A1(n18), .A2(n177), .ZN(tempResultB[123]) );
  NOR2_X1 U218 ( .A1(n22), .A2(n174), .ZN(tempResultB[153]) );
  NOR2_X1 U219 ( .A1(n16), .A2(n177), .ZN(tempResultB[124]) );
  NOR2_X1 U220 ( .A1(n24), .A2(n171), .ZN(tempResultB[184]) );
  NOR2_X1 U221 ( .A1(n14), .A2(n177), .ZN(tempResultB[125]) );
  NOR2_X1 U222 ( .A1(n18), .A2(n174), .ZN(tempResultB[155]) );
  NOR2_X1 U223 ( .A1(n22), .A2(n171), .ZN(tempResultB[185]) );
  NOR2_X1 U224 ( .A1(n16), .A2(n174), .ZN(tempResultB[156]) );
  NOR2_X1 U225 ( .A1(n20), .A2(n171), .ZN(tempResultB[186]) );
  NOR2_X1 U226 ( .A1(n14), .A2(n174), .ZN(tempResultB[157]) );
  NOR2_X1 U227 ( .A1(n18), .A2(n171), .ZN(tempResultB[187]) );
  NOR2_X1 U228 ( .A1(n16), .A2(n171), .ZN(tempResultB[188]) );
  NOR2_X1 U229 ( .A1(n14), .A2(n171), .ZN(tempResultB[189]) );
  NOR2_X1 U230 ( .A1(n39), .A2(n182), .ZN(tempResultB[50]) );
  NOR2_X1 U231 ( .A1(n27), .A2(n183), .ZN(tempResultB[55]) );
  NOR2_X1 U232 ( .A1(n86), .A2(n180), .ZN(tempResultB[66]) );
  NOR2_X1 U233 ( .A1(n41), .A2(n182), .ZN(tempResultB[49]) );
  NOR2_X1 U234 ( .A1(n44), .A2(n182), .ZN(tempResultB[48]) );
  NOR2_X1 U235 ( .A1(n33), .A2(n183), .ZN(tempResultB[52]) );
  NOR2_X1 U236 ( .A1(n56), .A2(n182), .ZN(tempResultB[44]) );
  NOR2_X1 U237 ( .A1(n53), .A2(n182), .ZN(tempResultB[45]) );
  NOR2_X1 U238 ( .A1(n47), .A2(n182), .ZN(tempResultB[47]) );
  NOR2_X1 U239 ( .A1(n50), .A2(n182), .ZN(tempResultB[46]) );
  NOR2_X1 U240 ( .A1(n36), .A2(n182), .ZN(tempResultB[51]) );
  NOR2_X1 U241 ( .A1(n62), .A2(n182), .ZN(tempResultB[42]) );
  NOR2_X1 U242 ( .A1(n89), .A2(n179), .ZN(tempResultB[65]) );
  NOR2_X1 U243 ( .A1(n90), .A2(n182), .ZN(tempResultB[33]) );
  NOR2_X1 U244 ( .A1(n87), .A2(n183), .ZN(tempResultB[34]) );
  NOR2_X1 U245 ( .A1(n21), .A2(n183), .ZN(tempResultB[58]) );
  NOR2_X1 U246 ( .A1(n89), .A2(n176), .ZN(tempResultB[97]) );
  NOR2_X1 U247 ( .A1(n86), .A2(n177), .ZN(tempResultB[98]) );
  NOR2_X1 U248 ( .A1(n89), .A2(n173), .ZN(tempResultB[129]) );
  NOR2_X1 U249 ( .A1(n86), .A2(n174), .ZN(tempResultB[130]) );
  NOR2_X1 U250 ( .A1(n89), .A2(n170), .ZN(tempResultB[161]) );
  NOR2_X1 U251 ( .A1(n86), .A2(n171), .ZN(tempResultB[162]) );
  NOR2_X1 U252 ( .A1(n89), .A2(n167), .ZN(tempResultB[193]) );
  NOR2_X1 U253 ( .A1(n86), .A2(n168), .ZN(tempResultB[194]) );
  NOR2_X1 U254 ( .A1(n61), .A2(n179), .ZN(tempResultB[74]) );
  NOR2_X1 U255 ( .A1(n89), .A2(n164), .ZN(tempResultB[225]) );
  NOR2_X1 U256 ( .A1(n86), .A2(n165), .ZN(tempResultB[226]) );
  NOR2_X1 U257 ( .A1(n61), .A2(n176), .ZN(tempResultB[106]) );
  NOR2_X1 U258 ( .A1(n55), .A2(n179), .ZN(tempResultB[76]) );
  NOR2_X1 U259 ( .A1(n89), .A2(n161), .ZN(tempResultB[257]) );
  NOR2_X1 U260 ( .A1(n52), .A2(n179), .ZN(tempResultB[77]) );
  NOR2_X1 U261 ( .A1(n61), .A2(n173), .ZN(tempResultB[138]) );
  NOR2_X1 U262 ( .A1(n55), .A2(n176), .ZN(tempResultB[108]) );
  NOR2_X1 U263 ( .A1(n49), .A2(n179), .ZN(tempResultB[78]) );
  NOR2_X1 U264 ( .A1(n52), .A2(n176), .ZN(tempResultB[109]) );
  NOR2_X1 U265 ( .A1(n46), .A2(n179), .ZN(tempResultB[79]) );
  NOR2_X1 U266 ( .A1(n61), .A2(n170), .ZN(tempResultB[170]) );
  NOR2_X1 U267 ( .A1(n55), .A2(n173), .ZN(tempResultB[140]) );
  NOR2_X1 U268 ( .A1(n49), .A2(n176), .ZN(tempResultB[110]) );
  NOR2_X1 U269 ( .A1(n43), .A2(n179), .ZN(tempResultB[80]) );
  NOR2_X1 U270 ( .A1(n52), .A2(n173), .ZN(tempResultB[141]) );
  NOR2_X1 U271 ( .A1(n46), .A2(n176), .ZN(tempResultB[111]) );
  NOR2_X1 U272 ( .A1(n40), .A2(n179), .ZN(tempResultB[81]) );
  NOR2_X1 U273 ( .A1(n55), .A2(n170), .ZN(tempResultB[172]) );
  NOR2_X1 U274 ( .A1(n49), .A2(n173), .ZN(tempResultB[142]) );
  NOR2_X1 U275 ( .A1(n43), .A2(n176), .ZN(tempResultB[112]) );
  NOR2_X1 U276 ( .A1(n52), .A2(n170), .ZN(tempResultB[173]) );
  NOR2_X1 U277 ( .A1(n46), .A2(n173), .ZN(tempResultB[143]) );
  NOR2_X1 U278 ( .A1(n40), .A2(n176), .ZN(tempResultB[113]) );
  NOR2_X1 U279 ( .A1(n35), .A2(n179), .ZN(tempResultB[83]) );
  NOR2_X1 U280 ( .A1(n49), .A2(n170), .ZN(tempResultB[174]) );
  NOR2_X1 U281 ( .A1(n43), .A2(n173), .ZN(tempResultB[144]) );
  NOR2_X1 U282 ( .A1(n46), .A2(n170), .ZN(tempResultB[175]) );
  NOR2_X1 U283 ( .A1(n40), .A2(n173), .ZN(tempResultB[145]) );
  NOR2_X1 U284 ( .A1(n35), .A2(n176), .ZN(tempResultB[115]) );
  NOR2_X1 U285 ( .A1(n43), .A2(n170), .ZN(tempResultB[176]) );
  NOR2_X1 U286 ( .A1(n40), .A2(n170), .ZN(tempResultB[177]) );
  NOR2_X1 U287 ( .A1(n35), .A2(n173), .ZN(tempResultB[147]) );
  NOR2_X1 U288 ( .A1(n35), .A2(n170), .ZN(tempResultB[179]) );
  NOR2_X1 U289 ( .A1(n17), .A2(n183), .ZN(tempResultB[60]) );
  NOR2_X1 U290 ( .A1(n38), .A2(n164), .ZN(tempResultB[242]) );
  NOR2_X1 U291 ( .A1(n26), .A2(n165), .ZN(tempResultB[247]) );
  NOR2_X1 U292 ( .A1(n26), .A2(n162), .ZN(tempResultB[279]) );
  NOR2_X1 U293 ( .A1(n32), .A2(n168), .ZN(tempResultB[212]) );
  NOR2_X1 U294 ( .A1(n32), .A2(n165), .ZN(tempResultB[244]) );
  NOR2_X1 U295 ( .A1(n159), .A2(n38), .ZN(tempResultB[306]) );
  NOR2_X1 U296 ( .A1(n159), .A2(n26), .ZN(tempResultB[311]) );
  NOR2_X1 U297 ( .A1(n159), .A2(n32), .ZN(tempResultB[308]) );
  NOR2_X1 U298 ( .A1(n160), .A2(n92), .ZN(tempResultB[288]) );
  NOR2_X1 U299 ( .A1(n94), .A2(n155), .ZN(tempResultB[320]) );
  NOR2_X1 U300 ( .A1(n94), .A2(n152), .ZN(tempResultB[352]) );
  NOR2_X1 U301 ( .A1(n94), .A2(n149), .ZN(tempResultB[384]) );
  NOR2_X1 U302 ( .A1(n94), .A2(n146), .ZN(tempResultB[416]) );
  NOR2_X1 U303 ( .A1(n94), .A2(n143), .ZN(tempResultB[448]) );
  NOR2_X1 U304 ( .A1(n94), .A2(n140), .ZN(tempResultB[480]) );
  NOR2_X1 U305 ( .A1(n12), .A2(n168), .ZN(tempResultB[222]) );
  NOR2_X1 U306 ( .A1(n12), .A2(n165), .ZN(tempResultB[254]) );
  NOR2_X1 U307 ( .A1(n12), .A2(n162), .ZN(tempResultB[286]) );
  NOR2_X1 U308 ( .A1(n9), .A2(n169), .ZN(tempResultB[223]) );
  NOR2_X1 U309 ( .A1(n9), .A2(n166), .ZN(tempResultB[255]) );
  NOR2_X1 U310 ( .A1(n9), .A2(n163), .ZN(tempResultB[287]) );
  NOR2_X1 U311 ( .A1(n158), .A2(n9), .ZN(tempResultB[319]) );
  NOR2_X1 U312 ( .A1(n58), .A2(n167), .ZN(tempResultB[203]) );
  NOR2_X1 U313 ( .A1(n58), .A2(n164), .ZN(tempResultB[235]) );
  NOR2_X1 U314 ( .A1(n58), .A2(n161), .ZN(tempResultB[267]) );
  NOR2_X1 U315 ( .A1(n91), .A2(n155), .ZN(tempResultB[321]) );
  NOR2_X1 U316 ( .A1(n91), .A2(n152), .ZN(tempResultB[353]) );
  NOR2_X1 U317 ( .A1(n91), .A2(n149), .ZN(tempResultB[385]) );
  NOR2_X1 U318 ( .A1(n91), .A2(n146), .ZN(tempResultB[417]) );
  NOR2_X1 U319 ( .A1(n160), .A2(n61), .ZN(tempResultB[298]) );
  NOR2_X1 U320 ( .A1(n91), .A2(n143), .ZN(tempResultB[449]) );
  NOR2_X1 U321 ( .A1(n160), .A2(n58), .ZN(tempResultB[299]) );
  NOR2_X1 U322 ( .A1(n160), .A2(n55), .ZN(tempResultB[300]) );
  NOR2_X1 U323 ( .A1(n91), .A2(n140), .ZN(tempResultB[481]) );
  NOR2_X1 U324 ( .A1(n160), .A2(n52), .ZN(tempResultB[301]) );
  NOR2_X1 U325 ( .A1(n160), .A2(n49), .ZN(tempResultB[302]) );
  NOR2_X1 U326 ( .A1(n160), .A2(n46), .ZN(tempResultB[303]) );
  NOR2_X1 U327 ( .A1(n160), .A2(n43), .ZN(tempResultB[304]) );
  NOR2_X1 U328 ( .A1(n158), .A2(n12), .ZN(tempResultB[318]) );
  NOR2_X1 U329 ( .A1(n74), .A2(n169), .ZN(tempResultB[198]) );
  NOR2_X1 U330 ( .A1(n80), .A2(n166), .ZN(tempResultB[228]) );
  NOR2_X1 U331 ( .A1(n71), .A2(n169), .ZN(tempResultB[199]) );
  NOR2_X1 U332 ( .A1(n77), .A2(n166), .ZN(tempResultB[229]) );
  NOR2_X1 U333 ( .A1(n83), .A2(n163), .ZN(tempResultB[259]) );
  NOR2_X1 U334 ( .A1(n67), .A2(n169), .ZN(tempResultB[200]) );
  NOR2_X1 U335 ( .A1(n74), .A2(n166), .ZN(tempResultB[230]) );
  NOR2_X1 U336 ( .A1(n80), .A2(n163), .ZN(tempResultB[260]) );
  NOR2_X1 U337 ( .A1(n71), .A2(n166), .ZN(tempResultB[231]) );
  NOR2_X1 U338 ( .A1(n77), .A2(n163), .ZN(tempResultB[261]) );
  NOR2_X1 U339 ( .A1(n64), .A2(n169), .ZN(tempResultB[201]) );
  NOR2_X1 U340 ( .A1(n67), .A2(n166), .ZN(tempResultB[232]) );
  NOR2_X1 U341 ( .A1(n74), .A2(n163), .ZN(tempResultB[262]) );
  NOR2_X1 U342 ( .A1(n71), .A2(n163), .ZN(tempResultB[263]) );
  NOR2_X1 U343 ( .A1(n64), .A2(n166), .ZN(tempResultB[233]) );
  NOR2_X1 U344 ( .A1(n67), .A2(n163), .ZN(tempResultB[264]) );
  NOR2_X1 U345 ( .A1(n64), .A2(n163), .ZN(tempResultB[265]) );
  NOR2_X1 U346 ( .A1(n30), .A2(n168), .ZN(tempResultB[213]) );
  NOR2_X1 U347 ( .A1(n30), .A2(n165), .ZN(tempResultB[245]) );
  NOR2_X1 U348 ( .A1(n24), .A2(n168), .ZN(tempResultB[216]) );
  NOR2_X1 U349 ( .A1(n28), .A2(n165), .ZN(tempResultB[246]) );
  NOR2_X1 U350 ( .A1(n22), .A2(n168), .ZN(tempResultB[217]) );
  NOR2_X1 U351 ( .A1(n30), .A2(n162), .ZN(tempResultB[277]) );
  NOR2_X1 U352 ( .A1(n20), .A2(n168), .ZN(tempResultB[218]) );
  NOR2_X1 U353 ( .A1(n24), .A2(n165), .ZN(tempResultB[248]) );
  NOR2_X1 U354 ( .A1(n18), .A2(n168), .ZN(tempResultB[219]) );
  NOR2_X1 U355 ( .A1(n22), .A2(n165), .ZN(tempResultB[249]) );
  NOR2_X1 U356 ( .A1(n16), .A2(n168), .ZN(tempResultB[220]) );
  NOR2_X1 U357 ( .A1(n20), .A2(n165), .ZN(tempResultB[250]) );
  NOR2_X1 U358 ( .A1(n24), .A2(n162), .ZN(tempResultB[280]) );
  NOR2_X1 U359 ( .A1(n14), .A2(n168), .ZN(tempResultB[221]) );
  NOR2_X1 U360 ( .A1(n18), .A2(n165), .ZN(tempResultB[251]) );
  NOR2_X1 U361 ( .A1(n22), .A2(n162), .ZN(tempResultB[281]) );
  NOR2_X1 U362 ( .A1(n16), .A2(n165), .ZN(tempResultB[252]) );
  NOR2_X1 U363 ( .A1(n20), .A2(n162), .ZN(tempResultB[282]) );
  NOR2_X1 U364 ( .A1(n14), .A2(n165), .ZN(tempResultB[253]) );
  NOR2_X1 U365 ( .A1(n18), .A2(n162), .ZN(tempResultB[283]) );
  NOR2_X1 U366 ( .A1(n16), .A2(n162), .ZN(tempResultB[284]) );
  NOR2_X1 U367 ( .A1(n14), .A2(n162), .ZN(tempResultB[285]) );
  NOR2_X1 U368 ( .A1(n159), .A2(n30), .ZN(tempResultB[309]) );
  NOR2_X1 U369 ( .A1(n159), .A2(n28), .ZN(tempResultB[310]) );
  NOR2_X1 U370 ( .A1(n159), .A2(n24), .ZN(tempResultB[312]) );
  NOR2_X1 U371 ( .A1(n159), .A2(n22), .ZN(tempResultB[313]) );
  NOR2_X1 U372 ( .A1(n159), .A2(n20), .ZN(tempResultB[314]) );
  NOR2_X1 U373 ( .A1(n159), .A2(n18), .ZN(tempResultB[315]) );
  NOR2_X1 U374 ( .A1(n158), .A2(n16), .ZN(tempResultB[316]) );
  NOR2_X1 U375 ( .A1(n158), .A2(n14), .ZN(tempResultB[317]) );
  NOR2_X1 U376 ( .A1(n86), .A2(n162), .ZN(tempResultB[258]) );
  NOR2_X1 U377 ( .A1(n159), .A2(n89), .ZN(tempResultB[289]) );
  NOR2_X1 U378 ( .A1(n158), .A2(n86), .ZN(tempResultB[290]) );
  NOR2_X1 U379 ( .A1(n158), .A2(n83), .ZN(tempResultB[291]) );
  NOR2_X1 U380 ( .A1(n158), .A2(n80), .ZN(tempResultB[292]) );
  NOR2_X1 U381 ( .A1(n61), .A2(n167), .ZN(tempResultB[202]) );
  NOR2_X1 U382 ( .A1(n158), .A2(n77), .ZN(tempResultB[293]) );
  NOR2_X1 U383 ( .A1(n158), .A2(n74), .ZN(tempResultB[294]) );
  NOR2_X1 U384 ( .A1(n61), .A2(n164), .ZN(tempResultB[234]) );
  NOR2_X1 U385 ( .A1(n55), .A2(n167), .ZN(tempResultB[204]) );
  NOR2_X1 U386 ( .A1(n158), .A2(n71), .ZN(tempResultB[295]) );
  NOR2_X1 U387 ( .A1(n52), .A2(n167), .ZN(tempResultB[205]) );
  NOR2_X1 U388 ( .A1(n158), .A2(n67), .ZN(tempResultB[296]) );
  NOR2_X1 U389 ( .A1(n61), .A2(n161), .ZN(tempResultB[266]) );
  NOR2_X1 U390 ( .A1(n55), .A2(n164), .ZN(tempResultB[236]) );
  NOR2_X1 U391 ( .A1(n49), .A2(n167), .ZN(tempResultB[206]) );
  NOR2_X1 U392 ( .A1(n64), .A2(n158), .ZN(tempResultB[297]) );
  NOR2_X1 U393 ( .A1(n52), .A2(n164), .ZN(tempResultB[237]) );
  NOR2_X1 U394 ( .A1(n46), .A2(n167), .ZN(tempResultB[207]) );
  NOR2_X1 U395 ( .A1(n55), .A2(n161), .ZN(tempResultB[268]) );
  NOR2_X1 U396 ( .A1(n49), .A2(n164), .ZN(tempResultB[238]) );
  NOR2_X1 U397 ( .A1(n43), .A2(n167), .ZN(tempResultB[208]) );
  NOR2_X1 U398 ( .A1(n52), .A2(n161), .ZN(tempResultB[269]) );
  NOR2_X1 U399 ( .A1(n46), .A2(n164), .ZN(tempResultB[239]) );
  NOR2_X1 U400 ( .A1(n40), .A2(n167), .ZN(tempResultB[209]) );
  NOR2_X1 U401 ( .A1(n49), .A2(n161), .ZN(tempResultB[270]) );
  NOR2_X1 U402 ( .A1(n43), .A2(n164), .ZN(tempResultB[240]) );
  NOR2_X1 U403 ( .A1(n46), .A2(n161), .ZN(tempResultB[271]) );
  NOR2_X1 U404 ( .A1(n40), .A2(n164), .ZN(tempResultB[241]) );
  NOR2_X1 U405 ( .A1(n35), .A2(n167), .ZN(tempResultB[211]) );
  NOR2_X1 U406 ( .A1(n43), .A2(n161), .ZN(tempResultB[272]) );
  NOR2_X1 U407 ( .A1(n35), .A2(n164), .ZN(tempResultB[243]) );
  NOR2_X1 U408 ( .A1(n40), .A2(n161), .ZN(tempResultB[273]) );
  NOR2_X1 U409 ( .A1(n35), .A2(n161), .ZN(tempResultB[275]) );
  NOR2_X1 U410 ( .A1(n159), .A2(n40), .ZN(tempResultB[305]) );
  NOR2_X1 U411 ( .A1(n159), .A2(n35), .ZN(tempResultB[307]) );
  NOR2_X1 U412 ( .A1(n11), .A2(n157), .ZN(tempResultB[351]) );
  NOR2_X1 U413 ( .A1(n11), .A2(n154), .ZN(tempResultB[383]) );
  NOR2_X1 U414 ( .A1(n11), .A2(n151), .ZN(tempResultB[415]) );
  NOR2_X1 U415 ( .A1(n11), .A2(n148), .ZN(tempResultB[447]) );
  NOR2_X1 U416 ( .A1(n11), .A2(n145), .ZN(tempResultB[479]) );
  NOR2_X1 U417 ( .A1(n93), .A2(n137), .ZN(tempResultB[512]) );
  NOR2_X1 U418 ( .A1(n93), .A2(n134), .ZN(tempResultB[544]) );
  NOR2_X1 U419 ( .A1(n93), .A2(n131), .ZN(tempResultB[576]) );
  NOR2_X1 U420 ( .A1(n93), .A2(n128), .ZN(tempResultB[608]) );
  NOR2_X1 U421 ( .A1(n93), .A2(n125), .ZN(tempResultB[640]) );
  NOR2_X1 U422 ( .A1(n93), .A2(n122), .ZN(tempResultB[672]) );
  NOR2_X1 U423 ( .A1(n84), .A2(n139), .ZN(tempResultB[515]) );
  NOR2_X1 U424 ( .A1(n81), .A2(n139), .ZN(tempResultB[516]) );
  NOR2_X1 U425 ( .A1(n78), .A2(n139), .ZN(tempResultB[517]) );
  NOR2_X1 U426 ( .A1(n84), .A2(n136), .ZN(tempResultB[547]) );
  NOR2_X1 U427 ( .A1(n75), .A2(n139), .ZN(tempResultB[518]) );
  NOR2_X1 U428 ( .A1(n81), .A2(n136), .ZN(tempResultB[548]) );
  NOR2_X1 U429 ( .A1(n72), .A2(n139), .ZN(tempResultB[519]) );
  NOR2_X1 U430 ( .A1(n78), .A2(n136), .ZN(tempResultB[549]) );
  NOR2_X1 U431 ( .A1(n84), .A2(n133), .ZN(tempResultB[579]) );
  NOR2_X1 U432 ( .A1(n69), .A2(n139), .ZN(tempResultB[520]) );
  NOR2_X1 U433 ( .A1(n75), .A2(n136), .ZN(tempResultB[550]) );
  NOR2_X1 U434 ( .A1(n81), .A2(n133), .ZN(tempResultB[580]) );
  NOR2_X1 U435 ( .A1(n72), .A2(n136), .ZN(tempResultB[551]) );
  NOR2_X1 U436 ( .A1(n78), .A2(n133), .ZN(tempResultB[581]) );
  NOR2_X1 U437 ( .A1(n84), .A2(n130), .ZN(tempResultB[611]) );
  NOR2_X1 U438 ( .A1(n65), .A2(n139), .ZN(tempResultB[521]) );
  NOR2_X1 U439 ( .A1(n69), .A2(n136), .ZN(tempResultB[552]) );
  NOR2_X1 U440 ( .A1(n75), .A2(n133), .ZN(tempResultB[582]) );
  NOR2_X1 U441 ( .A1(n81), .A2(n130), .ZN(tempResultB[612]) );
  NOR2_X1 U442 ( .A1(n72), .A2(n133), .ZN(tempResultB[583]) );
  NOR2_X1 U443 ( .A1(n84), .A2(n127), .ZN(tempResultB[643]) );
  NOR2_X1 U444 ( .A1(n65), .A2(n136), .ZN(tempResultB[553]) );
  NOR2_X1 U445 ( .A1(n69), .A2(n133), .ZN(tempResultB[584]) );
  NOR2_X1 U446 ( .A1(n75), .A2(n130), .ZN(tempResultB[614]) );
  NOR2_X1 U447 ( .A1(n81), .A2(n127), .ZN(tempResultB[644]) );
  NOR2_X1 U448 ( .A1(n90), .A2(n137), .ZN(tempResultB[513]) );
  NOR2_X1 U449 ( .A1(n87), .A2(n138), .ZN(tempResultB[514]) );
  NOR2_X1 U450 ( .A1(n90), .A2(n134), .ZN(tempResultB[545]) );
  NOR2_X1 U451 ( .A1(n87), .A2(n135), .ZN(tempResultB[546]) );
  NOR2_X1 U452 ( .A1(n90), .A2(n131), .ZN(tempResultB[577]) );
  NOR2_X1 U453 ( .A1(n87), .A2(n132), .ZN(tempResultB[578]) );
  NOR2_X1 U454 ( .A1(n90), .A2(n128), .ZN(tempResultB[609]) );
  NOR2_X1 U455 ( .A1(n87), .A2(n129), .ZN(tempResultB[610]) );
  NOR2_X1 U456 ( .A1(n90), .A2(n125), .ZN(tempResultB[641]) );
  NOR2_X1 U457 ( .A1(n87), .A2(n126), .ZN(tempResultB[642]) );
  NOR2_X1 U458 ( .A1(n62), .A2(n137), .ZN(tempResultB[522]) );
  NOR2_X1 U459 ( .A1(n90), .A2(n122), .ZN(tempResultB[673]) );
  NOR2_X1 U460 ( .A1(n87), .A2(n123), .ZN(tempResultB[674]) );
  NOR2_X1 U461 ( .A1(n62), .A2(n134), .ZN(tempResultB[554]) );
  NOR2_X1 U462 ( .A1(n56), .A2(n137), .ZN(tempResultB[524]) );
  NOR2_X1 U463 ( .A1(n31), .A2(n138), .ZN(tempResultB[533]) );
  NOR2_X1 U464 ( .A1(n31), .A2(n135), .ZN(tempResultB[565]) );
  NOR2_X1 U465 ( .A1(n31), .A2(n132), .ZN(tempResultB[597]) );
  NOR2_X1 U466 ( .A1(n31), .A2(n129), .ZN(tempResultB[629]) );
  NOR2_X1 U467 ( .A1(n15), .A2(n138), .ZN(tempResultB[541]) );
  NOR2_X1 U468 ( .A1(n29), .A2(n138), .ZN(tempResultB[534]) );
  NOR2_X1 U469 ( .A1(n29), .A2(n135), .ZN(tempResultB[566]) );
  NOR2_X1 U470 ( .A1(n23), .A2(n138), .ZN(tempResultB[537]) );
  NOR2_X1 U471 ( .A1(n29), .A2(n132), .ZN(tempResultB[598]) );
  NOR2_X1 U472 ( .A1(n19), .A2(n138), .ZN(tempResultB[539]) );
  NOR2_X1 U473 ( .A1(n23), .A2(n135), .ZN(tempResultB[569]) );
  NOR2_X1 U474 ( .A1(n19), .A2(n135), .ZN(tempResultB[571]) );
  NOR2_X1 U475 ( .A1(n23), .A2(n132), .ZN(tempResultB[601]) );
  NOR2_X1 U476 ( .A1(n15), .A2(n135), .ZN(tempResultB[573]) );
  NOR2_X1 U477 ( .A1(n19), .A2(n132), .ZN(tempResultB[603]) );
  NOR2_X1 U478 ( .A1(n15), .A2(n132), .ZN(tempResultB[605]) );
  NOR2_X1 U479 ( .A1(n11), .A2(n142), .ZN(tempResultB[511]) );
  NOR2_X1 U480 ( .A1(n13), .A2(n135), .ZN(tempResultB[574]) );
  NOR2_X1 U481 ( .A1(n13), .A2(n132), .ZN(tempResultB[606]) );
  NOR2_X1 U482 ( .A1(n10), .A2(n139), .ZN(tempResultB[543]) );
  NOR2_X1 U483 ( .A1(n10), .A2(n136), .ZN(tempResultB[575]) );
  NOR2_X1 U484 ( .A1(n10), .A2(n133), .ZN(tempResultB[607]) );
  NOR2_X1 U485 ( .A1(n93), .A2(n119), .ZN(tempResultB[704]) );
  NOR2_X1 U486 ( .A1(n93), .A2(n116), .ZN(tempResultB[736]) );
  NOR2_X1 U487 ( .A1(n93), .A2(n113), .ZN(tempResultB[768]) );
  NOR2_X1 U488 ( .A1(n93), .A2(n110), .ZN(tempResultB[800]) );
  NOR2_X1 U489 ( .A1(n93), .A2(n107), .ZN(tempResultB[832]) );
  NOR2_X1 U490 ( .A1(n92), .A2(n104), .ZN(tempResultB[864]) );
  NOR2_X1 U491 ( .A1(n92), .A2(n101), .ZN(tempResultB[896]) );
  NOR2_X1 U492 ( .A1(n59), .A2(n128), .ZN(tempResultB[619]) );
  NOR2_X1 U493 ( .A1(n59), .A2(n125), .ZN(tempResultB[651]) );
  NOR2_X1 U494 ( .A1(n59), .A2(n122), .ZN(tempResultB[683]) );
  NOR2_X1 U495 ( .A1(n59), .A2(n119), .ZN(tempResultB[715]) );
  NOR2_X1 U496 ( .A1(n25), .A2(n138), .ZN(tempResultB[536]) );
  NOR2_X1 U497 ( .A1(n59), .A2(n116), .ZN(tempResultB[747]) );
  NOR2_X1 U498 ( .A1(n25), .A2(n135), .ZN(tempResultB[568]) );
  NOR2_X1 U499 ( .A1(n25), .A2(n132), .ZN(tempResultB[600]) );
  NOR2_X1 U500 ( .A1(n13), .A2(n138), .ZN(tempResultB[542]) );
  NOR2_X1 U501 ( .A1(n72), .A2(n130), .ZN(tempResultB[615]) );
  NOR2_X1 U502 ( .A1(n78), .A2(n127), .ZN(tempResultB[645]) );
  NOR2_X1 U503 ( .A1(n84), .A2(n124), .ZN(tempResultB[675]) );
  NOR2_X1 U504 ( .A1(n69), .A2(n130), .ZN(tempResultB[616]) );
  NOR2_X1 U505 ( .A1(n75), .A2(n127), .ZN(tempResultB[646]) );
  NOR2_X1 U506 ( .A1(n81), .A2(n124), .ZN(tempResultB[676]) );
  NOR2_X1 U507 ( .A1(n72), .A2(n127), .ZN(tempResultB[647]) );
  NOR2_X1 U508 ( .A1(n78), .A2(n124), .ZN(tempResultB[677]) );
  NOR2_X1 U509 ( .A1(n84), .A2(n121), .ZN(tempResultB[707]) );
  NOR2_X1 U510 ( .A1(n65), .A2(n130), .ZN(tempResultB[617]) );
  NOR2_X1 U511 ( .A1(n69), .A2(n127), .ZN(tempResultB[648]) );
  NOR2_X1 U512 ( .A1(n75), .A2(n124), .ZN(tempResultB[678]) );
  NOR2_X1 U513 ( .A1(n81), .A2(n121), .ZN(tempResultB[708]) );
  NOR2_X1 U514 ( .A1(n72), .A2(n124), .ZN(tempResultB[679]) );
  NOR2_X1 U515 ( .A1(n78), .A2(n121), .ZN(tempResultB[709]) );
  NOR2_X1 U516 ( .A1(n84), .A2(n118), .ZN(tempResultB[739]) );
  NOR2_X1 U517 ( .A1(n69), .A2(n124), .ZN(tempResultB[680]) );
  NOR2_X1 U518 ( .A1(n75), .A2(n121), .ZN(tempResultB[710]) );
  NOR2_X1 U519 ( .A1(n81), .A2(n118), .ZN(tempResultB[740]) );
  NOR2_X1 U520 ( .A1(n72), .A2(n121), .ZN(tempResultB[711]) );
  NOR2_X1 U521 ( .A1(n78), .A2(n118), .ZN(tempResultB[741]) );
  NOR2_X1 U522 ( .A1(n84), .A2(n115), .ZN(tempResultB[771]) );
  NOR2_X1 U523 ( .A1(n65), .A2(n124), .ZN(tempResultB[681]) );
  NOR2_X1 U524 ( .A1(n69), .A2(n121), .ZN(tempResultB[712]) );
  NOR2_X1 U525 ( .A1(n75), .A2(n118), .ZN(tempResultB[742]) );
  NOR2_X1 U526 ( .A1(n81), .A2(n115), .ZN(tempResultB[772]) );
  NOR2_X1 U527 ( .A1(n72), .A2(n118), .ZN(tempResultB[743]) );
  NOR2_X1 U528 ( .A1(n78), .A2(n115), .ZN(tempResultB[773]) );
  NOR2_X1 U529 ( .A1(n84), .A2(n112), .ZN(tempResultB[803]) );
  NOR2_X1 U530 ( .A1(n65), .A2(n121), .ZN(tempResultB[713]) );
  NOR2_X1 U531 ( .A1(n69), .A2(n118), .ZN(tempResultB[744]) );
  NOR2_X1 U532 ( .A1(n75), .A2(n115), .ZN(tempResultB[774]) );
  NOR2_X1 U533 ( .A1(n81), .A2(n112), .ZN(tempResultB[804]) );
  NOR2_X1 U534 ( .A1(n78), .A2(n112), .ZN(tempResultB[805]) );
  NOR2_X1 U535 ( .A1(n84), .A2(n109), .ZN(tempResultB[835]) );
  NOR2_X1 U536 ( .A1(n65), .A2(n118), .ZN(tempResultB[745]) );
  NOR2_X1 U537 ( .A1(n69), .A2(n115), .ZN(tempResultB[776]) );
  NOR2_X1 U538 ( .A1(n75), .A2(n112), .ZN(tempResultB[806]) );
  NOR2_X1 U539 ( .A1(n81), .A2(n109), .ZN(tempResultB[836]) );
  NOR2_X1 U540 ( .A1(n72), .A2(n112), .ZN(tempResultB[807]) );
  NOR2_X1 U541 ( .A1(n78), .A2(n109), .ZN(tempResultB[837]) );
  NOR2_X1 U542 ( .A1(n83), .A2(n106), .ZN(tempResultB[867]) );
  NOR2_X1 U543 ( .A1(n65), .A2(n115), .ZN(tempResultB[777]) );
  NOR2_X1 U544 ( .A1(n69), .A2(n112), .ZN(tempResultB[808]) );
  NOR2_X1 U545 ( .A1(n75), .A2(n109), .ZN(tempResultB[838]) );
  NOR2_X1 U546 ( .A1(n80), .A2(n106), .ZN(tempResultB[868]) );
  NOR2_X1 U547 ( .A1(n39), .A2(n137), .ZN(tempResultB[530]) );
  NOR2_X1 U548 ( .A1(n39), .A2(n134), .ZN(tempResultB[562]) );
  NOR2_X1 U549 ( .A1(n39), .A2(n131), .ZN(tempResultB[594]) );
  NOR2_X1 U550 ( .A1(n27), .A2(n138), .ZN(tempResultB[535]) );
  NOR2_X1 U551 ( .A1(n39), .A2(n128), .ZN(tempResultB[626]) );
  NOR2_X1 U552 ( .A1(n27), .A2(n135), .ZN(tempResultB[567]) );
  NOR2_X1 U553 ( .A1(n27), .A2(n132), .ZN(tempResultB[599]) );
  NOR2_X1 U554 ( .A1(n90), .A2(n119), .ZN(tempResultB[705]) );
  NOR2_X1 U555 ( .A1(n53), .A2(n137), .ZN(tempResultB[525]) );
  NOR2_X1 U556 ( .A1(n87), .A2(n120), .ZN(tempResultB[706]) );
  NOR2_X1 U557 ( .A1(n50), .A2(n137), .ZN(tempResultB[526]) );
  NOR2_X1 U558 ( .A1(n62), .A2(n131), .ZN(tempResultB[586]) );
  NOR2_X1 U559 ( .A1(n56), .A2(n134), .ZN(tempResultB[556]) );
  NOR2_X1 U560 ( .A1(n90), .A2(n116), .ZN(tempResultB[737]) );
  NOR2_X1 U561 ( .A1(n47), .A2(n137), .ZN(tempResultB[527]) );
  NOR2_X1 U562 ( .A1(n53), .A2(n134), .ZN(tempResultB[557]) );
  NOR2_X1 U563 ( .A1(n87), .A2(n117), .ZN(tempResultB[738]) );
  NOR2_X1 U564 ( .A1(n44), .A2(n137), .ZN(tempResultB[528]) );
  NOR2_X1 U565 ( .A1(n62), .A2(n128), .ZN(tempResultB[618]) );
  NOR2_X1 U566 ( .A1(n50), .A2(n134), .ZN(tempResultB[558]) );
  NOR2_X1 U567 ( .A1(n56), .A2(n131), .ZN(tempResultB[588]) );
  NOR2_X1 U568 ( .A1(n90), .A2(n113), .ZN(tempResultB[769]) );
  NOR2_X1 U569 ( .A1(n41), .A2(n137), .ZN(tempResultB[529]) );
  NOR2_X1 U570 ( .A1(n47), .A2(n134), .ZN(tempResultB[559]) );
  NOR2_X1 U571 ( .A1(n53), .A2(n131), .ZN(tempResultB[589]) );
  NOR2_X1 U572 ( .A1(n87), .A2(n114), .ZN(tempResultB[770]) );
  NOR2_X1 U573 ( .A1(n44), .A2(n134), .ZN(tempResultB[560]) );
  NOR2_X1 U574 ( .A1(n50), .A2(n131), .ZN(tempResultB[590]) );
  NOR2_X1 U575 ( .A1(n56), .A2(n128), .ZN(tempResultB[620]) );
  NOR2_X1 U576 ( .A1(n62), .A2(n125), .ZN(tempResultB[650]) );
  NOR2_X1 U577 ( .A1(n90), .A2(n110), .ZN(tempResultB[801]) );
  NOR2_X1 U578 ( .A1(n36), .A2(n137), .ZN(tempResultB[531]) );
  NOR2_X1 U579 ( .A1(n41), .A2(n134), .ZN(tempResultB[561]) );
  NOR2_X1 U580 ( .A1(n47), .A2(n131), .ZN(tempResultB[591]) );
  NOR2_X1 U581 ( .A1(n53), .A2(n128), .ZN(tempResultB[621]) );
  NOR2_X1 U582 ( .A1(n87), .A2(n111), .ZN(tempResultB[802]) );
  NOR2_X1 U583 ( .A1(n33), .A2(n138), .ZN(tempResultB[532]) );
  NOR2_X1 U584 ( .A1(n44), .A2(n131), .ZN(tempResultB[592]) );
  NOR2_X1 U585 ( .A1(n50), .A2(n128), .ZN(tempResultB[622]) );
  NOR2_X1 U586 ( .A1(n56), .A2(n125), .ZN(tempResultB[652]) );
  NOR2_X1 U587 ( .A1(n62), .A2(n122), .ZN(tempResultB[682]) );
  NOR2_X1 U588 ( .A1(n90), .A2(n107), .ZN(tempResultB[833]) );
  NOR2_X1 U589 ( .A1(n36), .A2(n134), .ZN(tempResultB[563]) );
  NOR2_X1 U590 ( .A1(n41), .A2(n131), .ZN(tempResultB[593]) );
  NOR2_X1 U591 ( .A1(n47), .A2(n128), .ZN(tempResultB[623]) );
  NOR2_X1 U592 ( .A1(n53), .A2(n125), .ZN(tempResultB[653]) );
  NOR2_X1 U593 ( .A1(n87), .A2(n108), .ZN(tempResultB[834]) );
  NOR2_X1 U594 ( .A1(n33), .A2(n135), .ZN(tempResultB[564]) );
  NOR2_X1 U595 ( .A1(n44), .A2(n128), .ZN(tempResultB[624]) );
  NOR2_X1 U596 ( .A1(n50), .A2(n125), .ZN(tempResultB[654]) );
  NOR2_X1 U597 ( .A1(n56), .A2(n122), .ZN(tempResultB[684]) );
  NOR2_X1 U598 ( .A1(n62), .A2(n119), .ZN(tempResultB[714]) );
  NOR2_X1 U599 ( .A1(n89), .A2(n104), .ZN(tempResultB[865]) );
  NOR2_X1 U600 ( .A1(n36), .A2(n131), .ZN(tempResultB[595]) );
  NOR2_X1 U601 ( .A1(n41), .A2(n128), .ZN(tempResultB[625]) );
  NOR2_X1 U602 ( .A1(n47), .A2(n125), .ZN(tempResultB[655]) );
  NOR2_X1 U603 ( .A1(n53), .A2(n122), .ZN(tempResultB[685]) );
  NOR2_X1 U604 ( .A1(n86), .A2(n105), .ZN(tempResultB[866]) );
  NOR2_X1 U605 ( .A1(n33), .A2(n132), .ZN(tempResultB[596]) );
  NOR2_X1 U606 ( .A1(n44), .A2(n125), .ZN(tempResultB[656]) );
  NOR2_X1 U607 ( .A1(n50), .A2(n122), .ZN(tempResultB[686]) );
  NOR2_X1 U608 ( .A1(n56), .A2(n119), .ZN(tempResultB[716]) );
  NOR2_X1 U609 ( .A1(n62), .A2(n116), .ZN(tempResultB[746]) );
  NOR2_X1 U610 ( .A1(n89), .A2(n101), .ZN(tempResultB[897]) );
  NOR2_X1 U611 ( .A1(n36), .A2(n128), .ZN(tempResultB[627]) );
  NOR2_X1 U612 ( .A1(n41), .A2(n125), .ZN(tempResultB[657]) );
  NOR2_X1 U613 ( .A1(n47), .A2(n122), .ZN(tempResultB[687]) );
  NOR2_X1 U614 ( .A1(n53), .A2(n119), .ZN(tempResultB[717]) );
  NOR2_X1 U615 ( .A1(n86), .A2(n102), .ZN(tempResultB[898]) );
  NOR2_X1 U616 ( .A1(n21), .A2(n138), .ZN(tempResultB[538]) );
  NOR2_X1 U617 ( .A1(n56), .A2(n116), .ZN(tempResultB[748]) );
  NOR2_X1 U618 ( .A1(n62), .A2(n113), .ZN(tempResultB[778]) );
  NOR2_X1 U619 ( .A1(n17), .A2(n138), .ZN(tempResultB[540]) );
  NOR2_X1 U620 ( .A1(n21), .A2(n135), .ZN(tempResultB[570]) );
  NOR2_X1 U621 ( .A1(n17), .A2(n135), .ZN(tempResultB[572]) );
  NOR2_X1 U622 ( .A1(n21), .A2(n132), .ZN(tempResultB[602]) );
  NOR2_X1 U623 ( .A1(n17), .A2(n132), .ZN(tempResultB[604]) );
  NOR2_X1 U624 ( .A1(n31), .A2(n126), .ZN(tempResultB[661]) );
  NOR2_X1 U625 ( .A1(n31), .A2(n123), .ZN(tempResultB[693]) );
  NOR2_X1 U626 ( .A1(n31), .A2(n120), .ZN(tempResultB[725]) );
  NOR2_X1 U627 ( .A1(n31), .A2(n117), .ZN(tempResultB[757]) );
  NOR2_X1 U628 ( .A1(n31), .A2(n114), .ZN(tempResultB[789]) );
  NOR2_X1 U629 ( .A1(n31), .A2(n111), .ZN(tempResultB[821]) );
  BUF_X1 U630 ( .A(n192), .Z(n195) );
  NOR2_X1 U631 ( .A1(n29), .A2(n129), .ZN(tempResultB[630]) );
  NOR2_X1 U632 ( .A1(n29), .A2(n126), .ZN(tempResultB[662]) );
  NOR2_X1 U633 ( .A1(n23), .A2(n129), .ZN(tempResultB[633]) );
  NOR2_X1 U634 ( .A1(n29), .A2(n123), .ZN(tempResultB[694]) );
  NOR2_X1 U635 ( .A1(n19), .A2(n129), .ZN(tempResultB[635]) );
  NOR2_X1 U636 ( .A1(n23), .A2(n126), .ZN(tempResultB[665]) );
  NOR2_X1 U637 ( .A1(n29), .A2(n120), .ZN(tempResultB[726]) );
  NOR2_X1 U638 ( .A1(n15), .A2(n129), .ZN(tempResultB[637]) );
  NOR2_X1 U639 ( .A1(n19), .A2(n126), .ZN(tempResultB[667]) );
  NOR2_X1 U640 ( .A1(n23), .A2(n123), .ZN(tempResultB[697]) );
  NOR2_X1 U641 ( .A1(n29), .A2(n117), .ZN(tempResultB[758]) );
  NOR2_X1 U642 ( .A1(n15), .A2(n126), .ZN(tempResultB[669]) );
  NOR2_X1 U643 ( .A1(n19), .A2(n123), .ZN(tempResultB[699]) );
  NOR2_X1 U644 ( .A1(n23), .A2(n120), .ZN(tempResultB[729]) );
  NOR2_X1 U645 ( .A1(n29), .A2(n114), .ZN(tempResultB[790]) );
  NOR2_X1 U646 ( .A1(n15), .A2(n123), .ZN(tempResultB[701]) );
  NOR2_X1 U647 ( .A1(n19), .A2(n120), .ZN(tempResultB[731]) );
  NOR2_X1 U648 ( .A1(n23), .A2(n117), .ZN(tempResultB[761]) );
  NOR2_X1 U649 ( .A1(n15), .A2(n120), .ZN(tempResultB[733]) );
  NOR2_X1 U650 ( .A1(n19), .A2(n117), .ZN(tempResultB[763]) );
  NOR2_X1 U651 ( .A1(n15), .A2(n117), .ZN(tempResultB[765]) );
  NOR2_X1 U652 ( .A1(n13), .A2(n129), .ZN(tempResultB[638]) );
  NOR2_X1 U653 ( .A1(n13), .A2(n120), .ZN(tempResultB[734]) );
  NOR2_X1 U654 ( .A1(n13), .A2(n117), .ZN(tempResultB[766]) );
  NOR2_X1 U655 ( .A1(n10), .A2(n130), .ZN(tempResultB[639]) );
  NOR2_X1 U656 ( .A1(n10), .A2(n127), .ZN(tempResultB[671]) );
  NOR2_X1 U657 ( .A1(n10), .A2(n124), .ZN(tempResultB[703]) );
  NOR2_X1 U658 ( .A1(n10), .A2(n121), .ZN(tempResultB[735]) );
  NOR2_X1 U659 ( .A1(n92), .A2(n98), .ZN(tempResultB[928]) );
  NOR2_X1 U660 ( .A1(n58), .A2(n104), .ZN(tempResultB[875]) );
  NOR2_X1 U661 ( .A1(n58), .A2(n101), .ZN(tempResultB[907]) );
  NOR2_X1 U662 ( .A1(n58), .A2(n98), .ZN(tempResultB[939]) );
  NOR2_X1 U663 ( .A1(n59), .A2(n113), .ZN(tempResultB[779]) );
  NOR2_X1 U664 ( .A1(n59), .A2(n110), .ZN(tempResultB[811]) );
  NOR2_X1 U665 ( .A1(n25), .A2(n129), .ZN(tempResultB[632]) );
  NOR2_X1 U666 ( .A1(n59), .A2(n107), .ZN(tempResultB[843]) );
  NOR2_X1 U667 ( .A1(n25), .A2(n126), .ZN(tempResultB[664]) );
  NOR2_X1 U668 ( .A1(n25), .A2(n123), .ZN(tempResultB[696]) );
  NOR2_X1 U669 ( .A1(n25), .A2(n120), .ZN(tempResultB[728]) );
  NOR2_X1 U670 ( .A1(n13), .A2(n126), .ZN(tempResultB[670]) );
  NOR2_X1 U671 ( .A1(n25), .A2(n117), .ZN(tempResultB[760]) );
  NOR2_X1 U672 ( .A1(n13), .A2(n123), .ZN(tempResultB[702]) );
  NOR2_X1 U673 ( .A1(n72), .A2(n109), .ZN(tempResultB[839]) );
  NOR2_X1 U674 ( .A1(n77), .A2(n106), .ZN(tempResultB[869]) );
  NOR2_X1 U675 ( .A1(n65), .A2(n112), .ZN(tempResultB[809]) );
  NOR2_X1 U676 ( .A1(n69), .A2(n109), .ZN(tempResultB[840]) );
  NOR2_X1 U677 ( .A1(n74), .A2(n106), .ZN(tempResultB[870]) );
  NOR2_X1 U678 ( .A1(n80), .A2(n103), .ZN(tempResultB[900]) );
  NOR2_X1 U679 ( .A1(n71), .A2(n106), .ZN(tempResultB[871]) );
  NOR2_X1 U680 ( .A1(n77), .A2(n103), .ZN(tempResultB[901]) );
  NOR2_X1 U681 ( .A1(n83), .A2(n100), .ZN(tempResultB[931]) );
  NOR2_X1 U682 ( .A1(n65), .A2(n109), .ZN(tempResultB[841]) );
  NOR2_X1 U683 ( .A1(n67), .A2(n106), .ZN(tempResultB[872]) );
  NOR2_X1 U684 ( .A1(n74), .A2(n103), .ZN(tempResultB[902]) );
  NOR2_X1 U685 ( .A1(n80), .A2(n100), .ZN(tempResultB[932]) );
  NOR2_X1 U686 ( .A1(n71), .A2(n103), .ZN(tempResultB[903]) );
  NOR2_X1 U687 ( .A1(n83), .A2(n97), .ZN(tempResultB[963]) );
  NOR2_X1 U688 ( .A1(n64), .A2(n106), .ZN(tempResultB[873]) );
  NOR2_X1 U689 ( .A1(n74), .A2(n100), .ZN(tempResultB[934]) );
  NOR2_X1 U690 ( .A1(n80), .A2(n97), .ZN(tempResultB[964]) );
  NOR2_X1 U691 ( .A1(n71), .A2(n100), .ZN(tempResultB[935]) );
  NOR2_X1 U692 ( .A1(n77), .A2(n97), .ZN(tempResultB[965]) );
  NOR2_X1 U693 ( .A1(n64), .A2(n103), .ZN(tempResultB[905]) );
  NOR2_X1 U694 ( .A1(n67), .A2(n100), .ZN(tempResultB[936]) );
  NOR2_X1 U695 ( .A1(n74), .A2(n97), .ZN(tempResultB[966]) );
  NOR2_X1 U696 ( .A1(n71), .A2(n97), .ZN(tempResultB[967]) );
  NOR2_X1 U697 ( .A1(n64), .A2(n100), .ZN(tempResultB[937]) );
  NOR2_X1 U698 ( .A1(n67), .A2(n97), .ZN(tempResultB[968]) );
  NOR2_X1 U699 ( .A1(n64), .A2(n97), .ZN(tempResultB[969]) );
  NOR2_X1 U700 ( .A1(n39), .A2(n125), .ZN(tempResultB[658]) );
  NOR2_X1 U701 ( .A1(n39), .A2(n122), .ZN(tempResultB[690]) );
  NOR2_X1 U702 ( .A1(n27), .A2(n129), .ZN(tempResultB[631]) );
  NOR2_X1 U703 ( .A1(n39), .A2(n119), .ZN(tempResultB[722]) );
  NOR2_X1 U704 ( .A1(n27), .A2(n126), .ZN(tempResultB[663]) );
  NOR2_X1 U705 ( .A1(n39), .A2(n116), .ZN(tempResultB[754]) );
  NOR2_X1 U706 ( .A1(n27), .A2(n123), .ZN(tempResultB[695]) );
  NOR2_X1 U707 ( .A1(n39), .A2(n113), .ZN(tempResultB[786]) );
  NOR2_X1 U708 ( .A1(n27), .A2(n120), .ZN(tempResultB[727]) );
  NOR2_X1 U709 ( .A1(n39), .A2(n110), .ZN(tempResultB[818]) );
  NOR2_X1 U710 ( .A1(n27), .A2(n117), .ZN(tempResultB[759]) );
  NOR2_X1 U711 ( .A1(n39), .A2(n107), .ZN(tempResultB[850]) );
  NOR2_X1 U712 ( .A1(n33), .A2(n129), .ZN(tempResultB[628]) );
  NOR2_X1 U713 ( .A1(n44), .A2(n122), .ZN(tempResultB[688]) );
  NOR2_X1 U714 ( .A1(n50), .A2(n119), .ZN(tempResultB[718]) );
  NOR2_X1 U715 ( .A1(n89), .A2(n98), .ZN(tempResultB[929]) );
  NOR2_X1 U716 ( .A1(n36), .A2(n125), .ZN(tempResultB[659]) );
  NOR2_X1 U717 ( .A1(n41), .A2(n122), .ZN(tempResultB[689]) );
  NOR2_X1 U718 ( .A1(n47), .A2(n119), .ZN(tempResultB[719]) );
  NOR2_X1 U719 ( .A1(n53), .A2(n116), .ZN(tempResultB[749]) );
  NOR2_X1 U720 ( .A1(n86), .A2(n99), .ZN(tempResultB[930]) );
  NOR2_X1 U721 ( .A1(n92), .A2(n95), .ZN(tempResultB[960]) );
  NOR2_X1 U722 ( .A1(n33), .A2(n126), .ZN(tempResultB[660]) );
  NOR2_X1 U723 ( .A1(n44), .A2(n119), .ZN(tempResultB[720]) );
  NOR2_X1 U724 ( .A1(n50), .A2(n116), .ZN(tempResultB[750]) );
  NOR2_X1 U725 ( .A1(n56), .A2(n113), .ZN(tempResultB[780]) );
  NOR2_X1 U726 ( .A1(n62), .A2(n110), .ZN(tempResultB[810]) );
  NOR2_X1 U727 ( .A1(n89), .A2(n95), .ZN(tempResultB[961]) );
  NOR2_X1 U728 ( .A1(n36), .A2(n122), .ZN(tempResultB[691]) );
  NOR2_X1 U729 ( .A1(n41), .A2(n119), .ZN(tempResultB[721]) );
  NOR2_X1 U730 ( .A1(n47), .A2(n116), .ZN(tempResultB[751]) );
  NOR2_X1 U731 ( .A1(n53), .A2(n113), .ZN(tempResultB[781]) );
  NOR2_X1 U732 ( .A1(n86), .A2(n96), .ZN(tempResultB[962]) );
  NOR2_X1 U733 ( .A1(n33), .A2(n123), .ZN(tempResultB[692]) );
  NOR2_X1 U734 ( .A1(n44), .A2(n116), .ZN(tempResultB[752]) );
  NOR2_X1 U735 ( .A1(n50), .A2(n113), .ZN(tempResultB[782]) );
  NOR2_X1 U736 ( .A1(n56), .A2(n110), .ZN(tempResultB[812]) );
  NOR2_X1 U737 ( .A1(n62), .A2(n107), .ZN(tempResultB[842]) );
  NOR2_X1 U738 ( .A1(n36), .A2(n119), .ZN(tempResultB[723]) );
  NOR2_X1 U739 ( .A1(n41), .A2(n116), .ZN(tempResultB[753]) );
  NOR2_X1 U740 ( .A1(n47), .A2(n113), .ZN(tempResultB[783]) );
  NOR2_X1 U741 ( .A1(n53), .A2(n110), .ZN(tempResultB[813]) );
  NOR2_X1 U742 ( .A1(n21), .A2(n129), .ZN(tempResultB[634]) );
  NOR2_X1 U743 ( .A1(n44), .A2(n113), .ZN(tempResultB[784]) );
  NOR2_X1 U744 ( .A1(n50), .A2(n110), .ZN(tempResultB[814]) );
  NOR2_X1 U745 ( .A1(n56), .A2(n107), .ZN(tempResultB[844]) );
  NOR2_X1 U746 ( .A1(n61), .A2(n104), .ZN(tempResultB[874]) );
  NOR2_X1 U747 ( .A1(n36), .A2(n116), .ZN(tempResultB[755]) );
  NOR2_X1 U748 ( .A1(n53), .A2(n107), .ZN(tempResultB[845]) );
  NOR2_X1 U749 ( .A1(n17), .A2(n129), .ZN(tempResultB[636]) );
  NOR2_X1 U750 ( .A1(n21), .A2(n126), .ZN(tempResultB[666]) );
  NOR2_X1 U751 ( .A1(n33), .A2(n117), .ZN(tempResultB[756]) );
  NOR2_X1 U752 ( .A1(n44), .A2(n110), .ZN(tempResultB[816]) );
  NOR2_X1 U753 ( .A1(n50), .A2(n107), .ZN(tempResultB[846]) );
  NOR2_X1 U754 ( .A1(n61), .A2(n101), .ZN(tempResultB[906]) );
  NOR2_X1 U755 ( .A1(n36), .A2(n113), .ZN(tempResultB[787]) );
  NOR2_X1 U756 ( .A1(n41), .A2(n110), .ZN(tempResultB[817]) );
  NOR2_X1 U757 ( .A1(n17), .A2(n126), .ZN(tempResultB[668]) );
  NOR2_X1 U758 ( .A1(n21), .A2(n123), .ZN(tempResultB[698]) );
  NOR2_X1 U759 ( .A1(n49), .A2(n104), .ZN(tempResultB[878]) );
  NOR2_X1 U760 ( .A1(n47), .A2(n110), .ZN(tempResultB[815]) );
  NOR2_X1 U761 ( .A1(n55), .A2(n104), .ZN(tempResultB[876]) );
  NOR2_X1 U762 ( .A1(n47), .A2(n107), .ZN(tempResultB[847]) );
  NOR2_X1 U763 ( .A1(n52), .A2(n104), .ZN(tempResultB[877]) );
  NOR2_X1 U764 ( .A1(n33), .A2(n114), .ZN(tempResultB[788]) );
  NOR2_X1 U765 ( .A1(n44), .A2(n107), .ZN(tempResultB[848]) );
  NOR2_X1 U766 ( .A1(n55), .A2(n101), .ZN(tempResultB[908]) );
  NOR2_X1 U767 ( .A1(n61), .A2(n98), .ZN(tempResultB[938]) );
  NOR2_X1 U768 ( .A1(n36), .A2(n110), .ZN(tempResultB[819]) );
  NOR2_X1 U769 ( .A1(n41), .A2(n107), .ZN(tempResultB[849]) );
  NOR2_X1 U770 ( .A1(n46), .A2(n104), .ZN(tempResultB[879]) );
  NOR2_X1 U771 ( .A1(n52), .A2(n101), .ZN(tempResultB[909]) );
  NOR2_X1 U772 ( .A1(n61), .A2(n95), .ZN(tempResultB[970]) );
  NOR2_X1 U773 ( .A1(n21), .A2(n120), .ZN(tempResultB[730]) );
  NOR2_X1 U774 ( .A1(n43), .A2(n104), .ZN(tempResultB[880]) );
  NOR2_X1 U775 ( .A1(n49), .A2(n101), .ZN(tempResultB[910]) );
  NOR2_X1 U776 ( .A1(n33), .A2(n120), .ZN(tempResultB[724]) );
  NOR2_X1 U777 ( .A1(n41), .A2(n113), .ZN(tempResultB[785]) );
  NOR2_X1 U778 ( .A1(n17), .A2(n123), .ZN(tempResultB[700]) );
  NOR2_X1 U779 ( .A1(n33), .A2(n111), .ZN(tempResultB[820]) );
  NOR2_X1 U780 ( .A1(n55), .A2(n98), .ZN(tempResultB[940]) );
  NOR2_X1 U781 ( .A1(n36), .A2(n107), .ZN(tempResultB[851]) );
  NOR2_X1 U782 ( .A1(n40), .A2(n104), .ZN(tempResultB[881]) );
  NOR2_X1 U783 ( .A1(n52), .A2(n98), .ZN(tempResultB[941]) );
  NOR2_X1 U784 ( .A1(n17), .A2(n120), .ZN(tempResultB[732]) );
  NOR2_X1 U785 ( .A1(n21), .A2(n117), .ZN(tempResultB[762]) );
  NOR2_X1 U786 ( .A1(n17), .A2(n117), .ZN(tempResultB[764]) );
  NOR2_X1 U787 ( .A1(n38), .A2(n104), .ZN(tempResultB[882]) );
  NOR2_X1 U788 ( .A1(n38), .A2(n101), .ZN(tempResultB[914]) );
  NOR2_X1 U789 ( .A1(n38), .A2(n98), .ZN(tempResultB[946]) );
  NOR2_X1 U790 ( .A1(n26), .A2(n105), .ZN(tempResultB[887]) );
  NOR2_X1 U791 ( .A1(n38), .A2(n95), .ZN(tempResultB[978]) );
  NOR2_X1 U792 ( .A1(n26), .A2(n102), .ZN(tempResultB[919]) );
  NOR2_X1 U793 ( .A1(n26), .A2(n99), .ZN(tempResultB[951]) );
  NOR2_X1 U794 ( .A1(n32), .A2(n105), .ZN(tempResultB[884]) );
  NOR2_X1 U795 ( .A1(n32), .A2(n102), .ZN(tempResultB[916]) );
  NOR2_X1 U796 ( .A1(n32), .A2(n99), .ZN(tempResultB[948]) );
  NOR2_X1 U797 ( .A1(n32), .A2(n96), .ZN(tempResultB[980]) );
  NOR2_X1 U798 ( .A1(n31), .A2(n108), .ZN(tempResultB[853]) );
  BUF_X1 U799 ( .A(n192), .Z(n196) );
  NOR2_X1 U800 ( .A1(n29), .A2(n111), .ZN(tempResultB[822]) );
  NOR2_X1 U801 ( .A1(n23), .A2(n114), .ZN(tempResultB[793]) );
  NOR2_X1 U802 ( .A1(n29), .A2(n108), .ZN(tempResultB[854]) );
  NOR2_X1 U803 ( .A1(n19), .A2(n114), .ZN(tempResultB[795]) );
  NOR2_X1 U804 ( .A1(n23), .A2(n111), .ZN(tempResultB[825]) );
  NOR2_X1 U805 ( .A1(n15), .A2(n114), .ZN(tempResultB[797]) );
  NOR2_X1 U806 ( .A1(n19), .A2(n111), .ZN(tempResultB[827]) );
  NOR2_X1 U807 ( .A1(n23), .A2(n108), .ZN(tempResultB[857]) );
  NOR2_X1 U808 ( .A1(n15), .A2(n111), .ZN(tempResultB[829]) );
  NOR2_X1 U809 ( .A1(n19), .A2(n108), .ZN(tempResultB[859]) );
  NOR2_X1 U810 ( .A1(n15), .A2(n108), .ZN(tempResultB[861]) );
  NOR2_X1 U811 ( .A1(n12), .A2(n105), .ZN(tempResultB[894]) );
  NOR2_X1 U812 ( .A1(n10), .A2(n118), .ZN(tempResultB[767]) );
  NOR2_X1 U813 ( .A1(n10), .A2(n115), .ZN(tempResultB[799]) );
  NOR2_X1 U814 ( .A1(n10), .A2(n112), .ZN(tempResultB[831]) );
  NOR2_X1 U815 ( .A1(n10), .A2(n109), .ZN(tempResultB[863]) );
  NOR2_X1 U816 ( .A1(n18), .A2(n105), .ZN(tempResultB[891]) );
  NOR2_X1 U817 ( .A1(n16), .A2(n105), .ZN(tempResultB[892]) );
  NOR2_X1 U818 ( .A1(n17), .A2(n108), .ZN(tempResultB[860]) );
  NOR2_X1 U819 ( .A1(n58), .A2(n95), .ZN(tempResultB[971]) );
  NOR2_X1 U820 ( .A1(n25), .A2(n114), .ZN(tempResultB[792]) );
  NOR2_X1 U821 ( .A1(n25), .A2(n111), .ZN(tempResultB[824]) );
  NOR2_X1 U822 ( .A1(n25), .A2(n108), .ZN(tempResultB[856]) );
  NOR2_X1 U823 ( .A1(n13), .A2(n114), .ZN(tempResultB[798]) );
  NOR2_X1 U824 ( .A1(n13), .A2(n111), .ZN(tempResultB[830]) );
  NOR2_X1 U825 ( .A1(n13), .A2(n108), .ZN(tempResultB[862]) );
  NOR2_X1 U826 ( .A1(n30), .A2(n105), .ZN(tempResultB[885]) );
  NOR2_X1 U827 ( .A1(n28), .A2(n105), .ZN(tempResultB[886]) );
  NOR2_X1 U828 ( .A1(n30), .A2(n102), .ZN(tempResultB[917]) );
  NOR2_X1 U829 ( .A1(n24), .A2(n105), .ZN(tempResultB[888]) );
  NOR2_X1 U830 ( .A1(n28), .A2(n102), .ZN(tempResultB[918]) );
  NOR2_X1 U831 ( .A1(n22), .A2(n105), .ZN(tempResultB[889]) );
  NOR2_X1 U832 ( .A1(n30), .A2(n99), .ZN(tempResultB[949]) );
  NOR2_X1 U833 ( .A1(n20), .A2(n105), .ZN(tempResultB[890]) );
  NOR2_X1 U834 ( .A1(n24), .A2(n102), .ZN(tempResultB[920]) );
  NOR2_X1 U835 ( .A1(n28), .A2(n99), .ZN(tempResultB[950]) );
  NOR2_X1 U836 ( .A1(n22), .A2(n102), .ZN(tempResultB[921]) );
  NOR2_X1 U837 ( .A1(n30), .A2(n96), .ZN(tempResultB[981]) );
  NOR2_X1 U838 ( .A1(n20), .A2(n102), .ZN(tempResultB[922]) );
  NOR2_X1 U839 ( .A1(n24), .A2(n99), .ZN(tempResultB[952]) );
  NOR2_X1 U840 ( .A1(n28), .A2(n96), .ZN(tempResultB[982]) );
  NOR2_X1 U841 ( .A1(n14), .A2(n105), .ZN(tempResultB[893]) );
  NOR2_X1 U842 ( .A1(n18), .A2(n102), .ZN(tempResultB[923]) );
  NOR2_X1 U843 ( .A1(n22), .A2(n99), .ZN(tempResultB[953]) );
  NOR2_X1 U844 ( .A1(n27), .A2(n114), .ZN(tempResultB[791]) );
  NOR2_X1 U845 ( .A1(n27), .A2(n111), .ZN(tempResultB[823]) );
  NOR2_X1 U846 ( .A1(n27), .A2(n108), .ZN(tempResultB[855]) );
  NOR2_X1 U847 ( .A1(n46), .A2(n101), .ZN(tempResultB[911]) );
  NOR2_X1 U848 ( .A1(n55), .A2(n95), .ZN(tempResultB[972]) );
  NOR2_X1 U849 ( .A1(n43), .A2(n101), .ZN(tempResultB[912]) );
  NOR2_X1 U850 ( .A1(n49), .A2(n98), .ZN(tempResultB[942]) );
  NOR2_X1 U851 ( .A1(n52), .A2(n95), .ZN(tempResultB[973]) );
  NOR2_X1 U852 ( .A1(n35), .A2(n104), .ZN(tempResultB[883]) );
  NOR2_X1 U853 ( .A1(n40), .A2(n101), .ZN(tempResultB[913]) );
  NOR2_X1 U854 ( .A1(n49), .A2(n95), .ZN(tempResultB[974]) );
  NOR2_X1 U855 ( .A1(n33), .A2(n108), .ZN(tempResultB[852]) );
  NOR2_X1 U856 ( .A1(n46), .A2(n98), .ZN(tempResultB[943]) );
  NOR2_X1 U857 ( .A1(n21), .A2(n114), .ZN(tempResultB[794]) );
  NOR2_X1 U858 ( .A1(n43), .A2(n98), .ZN(tempResultB[944]) );
  NOR2_X1 U859 ( .A1(n46), .A2(n95), .ZN(tempResultB[975]) );
  NOR2_X1 U860 ( .A1(n35), .A2(n101), .ZN(tempResultB[915]) );
  NOR2_X1 U861 ( .A1(n40), .A2(n98), .ZN(tempResultB[945]) );
  NOR2_X1 U862 ( .A1(n43), .A2(n95), .ZN(tempResultB[976]) );
  NOR2_X1 U863 ( .A1(n21), .A2(n111), .ZN(tempResultB[826]) );
  NOR2_X1 U864 ( .A1(n40), .A2(n95), .ZN(tempResultB[977]) );
  NOR2_X1 U865 ( .A1(n35), .A2(n98), .ZN(tempResultB[947]) );
  NOR2_X1 U866 ( .A1(n35), .A2(n95), .ZN(tempResultB[979]) );
  NOR2_X1 U867 ( .A1(n17), .A2(n114), .ZN(tempResultB[796]) );
  NOR2_X1 U868 ( .A1(n17), .A2(n111), .ZN(tempResultB[828]) );
  NOR2_X1 U869 ( .A1(n21), .A2(n108), .ZN(tempResultB[858]) );
  NOR2_X1 U870 ( .A1(n26), .A2(n96), .ZN(tempResultB[983]) );
  NOR2_X1 U871 ( .A1(n12), .A2(n99), .ZN(tempResultB[958]) );
  NOR2_X1 U872 ( .A1(n12), .A2(n96), .ZN(tempResultB[990]) );
  NOR2_X1 U873 ( .A1(n12), .A2(n102), .ZN(tempResultB[926]) );
  NOR2_X1 U874 ( .A1(n9), .A2(n106), .ZN(tempResultB[895]) );
  NOR2_X1 U875 ( .A1(n9), .A2(n103), .ZN(tempResultB[927]) );
  NOR2_X1 U876 ( .A1(n9), .A2(n100), .ZN(tempResultB[959]) );
  NOR2_X1 U877 ( .A1(n9), .A2(n97), .ZN(tempResultB[991]) );
  NOR2_X1 U878 ( .A1(n16), .A2(n102), .ZN(tempResultB[924]) );
  NOR2_X1 U879 ( .A1(n20), .A2(n99), .ZN(tempResultB[954]) );
  NOR2_X1 U880 ( .A1(n24), .A2(n96), .ZN(tempResultB[984]) );
  NOR2_X1 U881 ( .A1(n14), .A2(n102), .ZN(tempResultB[925]) );
  NOR2_X1 U882 ( .A1(n18), .A2(n99), .ZN(tempResultB[955]) );
  NOR2_X1 U883 ( .A1(n22), .A2(n96), .ZN(tempResultB[985]) );
  NOR2_X1 U884 ( .A1(n16), .A2(n99), .ZN(tempResultB[956]) );
  NOR2_X1 U885 ( .A1(n20), .A2(n96), .ZN(tempResultB[986]) );
  NOR2_X1 U886 ( .A1(n14), .A2(n99), .ZN(tempResultB[957]) );
  NOR2_X1 U887 ( .A1(n18), .A2(n96), .ZN(tempResultB[987]) );
  NOR2_X1 U888 ( .A1(n16), .A2(n96), .ZN(tempResultB[988]) );
  NOR2_X1 U889 ( .A1(n14), .A2(n96), .ZN(tempResultB[989]) );
  BUF_X1 U890 ( .A(n191), .Z(n194) );
  BUF_X1 U891 ( .A(n220), .Z(n58) );
  BUF_X1 U892 ( .A(n207), .Z(n25) );
  BUF_X1 U893 ( .A(n210), .Z(n30) );
  BUF_X1 U894 ( .A(n259), .Z(n178) );
  BUF_X1 U895 ( .A(n258), .Z(n175) );
  BUF_X1 U896 ( .A(n257), .Z(n172) );
  BUF_X1 U897 ( .A(n256), .Z(n169) );
  BUF_X1 U898 ( .A(n255), .Z(n166) );
  BUF_X1 U899 ( .A(n230), .Z(n91) );
  BUF_X1 U900 ( .A(n231), .Z(n94) );
  BUF_X1 U901 ( .A(n258), .Z(n173) );
  BUF_X1 U902 ( .A(n257), .Z(n170) );
  BUF_X1 U903 ( .A(n256), .Z(n167) );
  BUF_X1 U904 ( .A(n255), .Z(n164) );
  BUF_X1 U905 ( .A(n254), .Z(n161) );
  BUF_X1 U906 ( .A(n259), .Z(n177) );
  BUF_X1 U907 ( .A(n258), .Z(n174) );
  BUF_X1 U908 ( .A(n257), .Z(n171) );
  BUF_X1 U909 ( .A(n256), .Z(n168) );
  BUF_X1 U910 ( .A(n255), .Z(n165) );
  CLKBUF_X1 U911 ( .A(n227), .Z(n80) );
  BUF_X1 U912 ( .A(n217), .Z(n49) );
  BUF_X1 U913 ( .A(n212), .Z(n35) );
  BUF_X1 U914 ( .A(n224), .Z(n71) );
  CLKBUF_X1 U915 ( .A(n231), .Z(n92) );
  CLKBUF_X1 U916 ( .A(n230), .Z(n89) );
  BUF_X1 U917 ( .A(n229), .Z(n86) );
  BUF_X1 U918 ( .A(n228), .Z(n83) );
  BUF_X1 U919 ( .A(n226), .Z(n77) );
  BUF_X1 U920 ( .A(n225), .Z(n74) );
  BUF_X1 U921 ( .A(n223), .Z(n67) );
  BUF_X1 U922 ( .A(n221), .Z(n61) );
  BUF_X1 U923 ( .A(n219), .Z(n55) );
  BUF_X1 U924 ( .A(n218), .Z(n52) );
  BUF_X1 U925 ( .A(n216), .Z(n46) );
  BUF_X1 U926 ( .A(n215), .Z(n43) );
  BUF_X1 U927 ( .A(n214), .Z(n40) );
  CLKBUF_X1 U928 ( .A(n200), .Z(n9) );
  BUF_X1 U929 ( .A(n205), .Z(n21) );
  BUF_X1 U930 ( .A(n222), .Z(n64) );
  BUF_X1 U931 ( .A(n203), .Z(n17) );
  BUF_X1 U932 ( .A(n263), .Z(n190) );
  BUF_X1 U933 ( .A(n212), .Z(n37) );
  BUF_X1 U934 ( .A(n217), .Z(n51) );
  BUF_X1 U935 ( .A(n211), .Z(n34) );
  BUF_X1 U936 ( .A(n220), .Z(n60) );
  BUF_X1 U937 ( .A(n216), .Z(n48) );
  BUF_X1 U938 ( .A(n222), .Z(n66) );
  BUF_X1 U939 ( .A(n224), .Z(n73) );
  BUF_X1 U940 ( .A(n214), .Z(n42) );
  BUF_X1 U941 ( .A(n215), .Z(n45) );
  BUF_X1 U942 ( .A(n221), .Z(n63) );
  BUF_X1 U943 ( .A(n219), .Z(n57) );
  BUF_X1 U944 ( .A(n226), .Z(n79) );
  BUF_X1 U945 ( .A(n228), .Z(n85) );
  BUF_X1 U946 ( .A(n223), .Z(n70) );
  BUF_X1 U947 ( .A(n225), .Z(n76) );
  BUF_X1 U948 ( .A(n229), .Z(n88) );
  BUF_X1 U949 ( .A(n263), .Z(n188) );
  BUF_X1 U950 ( .A(n263), .Z(n189) );
  BUF_X1 U951 ( .A(n262), .Z(n186) );
  BUF_X1 U952 ( .A(n254), .Z(n163) );
  BUF_X1 U953 ( .A(n253), .Z(n160) );
  BUF_X1 U954 ( .A(n254), .Z(n162) );
  BUF_X1 U955 ( .A(n253), .Z(n158) );
  BUF_X1 U956 ( .A(n253), .Z(n159) );
  BUF_X1 U957 ( .A(n252), .Z(n157) );
  BUF_X1 U958 ( .A(n251), .Z(n154) );
  BUF_X1 U959 ( .A(n250), .Z(n151) );
  BUF_X1 U960 ( .A(n249), .Z(n148) );
  BUF_X1 U961 ( .A(n252), .Z(n155) );
  BUF_X1 U962 ( .A(n251), .Z(n152) );
  BUF_X1 U963 ( .A(n250), .Z(n149) );
  BUF_X1 U964 ( .A(n249), .Z(n146) );
  BUF_X1 U965 ( .A(n248), .Z(n143) );
  BUF_X1 U966 ( .A(n247), .Z(n140) );
  BUF_X1 U967 ( .A(n252), .Z(n156) );
  BUF_X1 U968 ( .A(n251), .Z(n153) );
  BUF_X1 U969 ( .A(n250), .Z(n150) );
  BUF_X1 U970 ( .A(n249), .Z(n147) );
  BUF_X1 U971 ( .A(n248), .Z(n144) );
  BUF_X1 U972 ( .A(n246), .Z(n139) );
  BUF_X1 U973 ( .A(n245), .Z(n136) );
  BUF_X1 U974 ( .A(n244), .Z(n133) );
  BUF_X1 U975 ( .A(n243), .Z(n130) );
  BUF_X1 U976 ( .A(n242), .Z(n127) );
  BUF_X1 U977 ( .A(n246), .Z(n137) );
  BUF_X1 U978 ( .A(n245), .Z(n134) );
  BUF_X1 U979 ( .A(n244), .Z(n131) );
  BUF_X1 U980 ( .A(n243), .Z(n128) );
  BUF_X1 U981 ( .A(n242), .Z(n125) );
  BUF_X1 U982 ( .A(n241), .Z(n122) );
  BUF_X1 U983 ( .A(n246), .Z(n138) );
  BUF_X1 U984 ( .A(n245), .Z(n135) );
  BUF_X1 U985 ( .A(n244), .Z(n132) );
  BUF_X1 U986 ( .A(n243), .Z(n129) );
  BUF_X1 U987 ( .A(n242), .Z(n126) );
  BUF_X1 U988 ( .A(n241), .Z(n123) );
  BUF_X1 U989 ( .A(n248), .Z(n145) );
  BUF_X1 U990 ( .A(n247), .Z(n142) );
  BUF_X1 U991 ( .A(n247), .Z(n141) );
  BUF_X1 U992 ( .A(n241), .Z(n124) );
  BUF_X1 U993 ( .A(n240), .Z(n121) );
  BUF_X1 U994 ( .A(n239), .Z(n118) );
  BUF_X1 U995 ( .A(n238), .Z(n115) );
  BUF_X1 U996 ( .A(n237), .Z(n112) );
  BUF_X1 U997 ( .A(n236), .Z(n109) );
  BUF_X1 U998 ( .A(n235), .Z(n106) );
  BUF_X1 U999 ( .A(n234), .Z(n103) );
  BUF_X1 U1000 ( .A(n233), .Z(n100) );
  BUF_X1 U1001 ( .A(n240), .Z(n119) );
  BUF_X1 U1002 ( .A(n239), .Z(n116) );
  BUF_X1 U1003 ( .A(n238), .Z(n113) );
  BUF_X1 U1004 ( .A(n237), .Z(n110) );
  BUF_X1 U1005 ( .A(n236), .Z(n107) );
  BUF_X1 U1006 ( .A(n235), .Z(n104) );
  BUF_X1 U1007 ( .A(n234), .Z(n101) );
  BUF_X1 U1008 ( .A(n240), .Z(n120) );
  BUF_X1 U1009 ( .A(n239), .Z(n117) );
  BUF_X1 U1010 ( .A(n238), .Z(n114) );
  BUF_X1 U1011 ( .A(n237), .Z(n111) );
  BUF_X1 U1012 ( .A(n236), .Z(n108) );
  BUF_X1 U1013 ( .A(n235), .Z(n105) );
  BUF_X1 U1014 ( .A(n234), .Z(n102) );
  BUF_X1 U1015 ( .A(n232), .Z(n97) );
  BUF_X1 U1016 ( .A(n233), .Z(n98) );
  BUF_X1 U1017 ( .A(n232), .Z(n95) );
  BUF_X1 U1018 ( .A(n233), .Z(n99) );
  BUF_X1 U1019 ( .A(n232), .Z(n96) );
  INV_X1 U1020 ( .A(b_abs[0]), .ZN(n263) );
  INV_X1 U1021 ( .A(b_abs[1]), .ZN(n262) );
  NOR2_X1 U1022 ( .A1(n94), .A2(n188), .ZN(n68) );
  INV_X1 U1023 ( .A(a_abs[19]), .ZN(n212) );
  INV_X1 U1024 ( .A(a_abs[18]), .ZN(n213) );
  CLKBUF_X1 U1025 ( .A(n213), .Z(n38) );
  CLKBUF_X1 U1026 ( .A(n210), .Z(n31) );
  CLKBUF_X1 U1027 ( .A(n211), .Z(n32) );
  BUF_X1 U1028 ( .A(n209), .Z(n29) );
  INV_X1 U1029 ( .A(a_abs[22]), .ZN(n209) );
  BUF_X1 U1030 ( .A(n206), .Z(n23) );
  CLKBUF_X1 U1031 ( .A(n208), .Z(n26) );
  CLKBUF_X1 U1032 ( .A(n8), .Z(n4) );
  BUF_X2 U1033 ( .A(n8), .Z(n5) );
  BUF_X1 U1034 ( .A(a[31]), .Z(n8) );
  CLKBUF_X1 U1035 ( .A(a[31]), .Z(n199) );
  CLKBUF_X1 U1036 ( .A(n199), .Z(n6) );
  BUF_X2 U1037 ( .A(n199), .Z(n7) );
  BUF_X1 U1038 ( .A(n204), .Z(n19) );
  BUF_X1 U1039 ( .A(n202), .Z(n15) );
  NOR2_X1 U1040 ( .A1(n51), .A2(n140), .ZN(tempResultB[494]) );
  NOR2_X1 U1041 ( .A1(n51), .A2(n143), .ZN(tempResultB[462]) );
  NOR2_X1 U1042 ( .A1(n51), .A2(n146), .ZN(tempResultB[430]) );
  NOR2_X1 U1043 ( .A1(n51), .A2(n149), .ZN(tempResultB[398]) );
  NOR2_X1 U1044 ( .A1(n51), .A2(n152), .ZN(tempResultB[366]) );
  NOR2_X1 U1045 ( .A1(n51), .A2(n155), .ZN(tempResultB[334]) );
  NOR2_X1 U1046 ( .A1(n51), .A2(n185), .ZN(tempResultB[14]) );
  INV_X1 U1047 ( .A(a_abs[26]), .ZN(n205) );
  INV_X1 U1048 ( .A(a_abs[30]), .ZN(n201) );
  NOR2_X1 U1049 ( .A1(n30), .A2(n141), .ZN(tempResultB[501]) );
  NOR2_X1 U1050 ( .A1(n30), .A2(n144), .ZN(tempResultB[469]) );
  NOR2_X1 U1051 ( .A1(n30), .A2(n147), .ZN(tempResultB[437]) );
  NOR2_X1 U1052 ( .A1(n30), .A2(n150), .ZN(tempResultB[405]) );
  NOR2_X1 U1053 ( .A1(n30), .A2(n153), .ZN(tempResultB[373]) );
  NOR2_X1 U1054 ( .A1(n30), .A2(n156), .ZN(tempResultB[341]) );
  NOR2_X1 U1055 ( .A1(n210), .A2(n186), .ZN(tempResultB[21]) );
  NOR2_X1 U1056 ( .A1(n34), .A2(n141), .ZN(tempResultB[500]) );
  NOR2_X1 U1057 ( .A1(n34), .A2(n144), .ZN(tempResultB[468]) );
  NOR2_X1 U1058 ( .A1(n34), .A2(n147), .ZN(tempResultB[436]) );
  NOR2_X1 U1059 ( .A1(n34), .A2(n150), .ZN(tempResultB[404]) );
  NOR2_X1 U1060 ( .A1(n34), .A2(n153), .ZN(tempResultB[372]) );
  NOR2_X1 U1061 ( .A1(n34), .A2(n156), .ZN(tempResultB[340]) );
  NOR2_X1 U1062 ( .A1(n34), .A2(n186), .ZN(tempResultB[20]) );
  NOR2_X1 U1063 ( .A1(n34), .A2(n188), .ZN(tempResultA_0__19_) );
  INV_X1 U1064 ( .A(a_abs[29]), .ZN(n202) );
  NOR2_X1 U1065 ( .A1(n18), .A2(n141), .ZN(tempResultB[507]) );
  NOR2_X1 U1066 ( .A1(n18), .A2(n144), .ZN(tempResultB[475]) );
  NOR2_X1 U1067 ( .A1(n18), .A2(n147), .ZN(tempResultB[443]) );
  NOR2_X1 U1068 ( .A1(n18), .A2(n150), .ZN(tempResultB[411]) );
  NOR2_X1 U1069 ( .A1(n18), .A2(n153), .ZN(tempResultB[379]) );
  NOR2_X1 U1070 ( .A1(n18), .A2(n156), .ZN(tempResultB[347]) );
  NOR2_X1 U1071 ( .A1(n204), .A2(n186), .ZN(tempResultB[27]) );
  NOR2_X1 U1072 ( .A1(n63), .A2(n140), .ZN(tempResultB[490]) );
  NOR2_X1 U1073 ( .A1(n63), .A2(n143), .ZN(tempResultB[458]) );
  NOR2_X1 U1074 ( .A1(n63), .A2(n146), .ZN(tempResultB[426]) );
  NOR2_X1 U1075 ( .A1(n63), .A2(n149), .ZN(tempResultB[394]) );
  NOR2_X1 U1076 ( .A1(n63), .A2(n152), .ZN(tempResultB[362]) );
  NOR2_X1 U1077 ( .A1(n63), .A2(n155), .ZN(tempResultB[330]) );
  NOR2_X1 U1078 ( .A1(n63), .A2(n185), .ZN(tempResultB[10]) );
  NOR2_X1 U1079 ( .A1(n63), .A2(n190), .ZN(tempResultA_0__9_) );
  NOR2_X1 U1080 ( .A1(n37), .A2(n140), .ZN(tempResultB[499]) );
  NOR2_X1 U1081 ( .A1(n37), .A2(n143), .ZN(tempResultB[467]) );
  NOR2_X1 U1082 ( .A1(n37), .A2(n146), .ZN(tempResultB[435]) );
  NOR2_X1 U1083 ( .A1(n37), .A2(n149), .ZN(tempResultB[403]) );
  NOR2_X1 U1084 ( .A1(n37), .A2(n152), .ZN(tempResultB[371]) );
  NOR2_X1 U1085 ( .A1(n37), .A2(n155), .ZN(tempResultB[339]) );
  NOR2_X1 U1086 ( .A1(n37), .A2(n185), .ZN(tempResultB[19]) );
  NOR2_X1 U1087 ( .A1(n37), .A2(n188), .ZN(tempResultA_0__18_) );
  INV_X1 U1088 ( .A(a_abs[27]), .ZN(n204) );
  INV_X1 U1089 ( .A(a_abs[23]), .ZN(n208) );
  NOR2_X1 U1090 ( .A1(n14), .A2(n141), .ZN(tempResultB[509]) );
  NOR2_X1 U1091 ( .A1(n14), .A2(n144), .ZN(tempResultB[477]) );
  NOR2_X1 U1092 ( .A1(n14), .A2(n147), .ZN(tempResultB[445]) );
  NOR2_X1 U1101 ( .A1(n14), .A2(n150), .ZN(tempResultB[413]) );
  NOR2_X1 U1170 ( .A1(n14), .A2(n153), .ZN(tempResultB[381]) );
  NOR2_X1 U1220 ( .A1(n14), .A2(n156), .ZN(tempResultB[349]) );
  NOR2_X1 U1221 ( .A1(n202), .A2(n186), .ZN(tempResultB[29]) );
  NOR2_X1 U1222 ( .A1(n16), .A2(n141), .ZN(tempResultB[508]) );
  NOR2_X1 U1223 ( .A1(n16), .A2(n144), .ZN(tempResultB[476]) );
  NOR2_X1 U1224 ( .A1(n16), .A2(n147), .ZN(tempResultB[444]) );
  NOR2_X1 U1225 ( .A1(n16), .A2(n150), .ZN(tempResultB[412]) );
  NOR2_X1 U1226 ( .A1(n16), .A2(n153), .ZN(tempResultB[380]) );
  NOR2_X1 U1227 ( .A1(n16), .A2(n156), .ZN(tempResultB[348]) );
  NOR2_X1 U1228 ( .A1(n203), .A2(n186), .ZN(tempResultB[28]) );
  INV_X1 U1229 ( .A(a_abs[24]), .ZN(n207) );
  NOR2_X1 U1230 ( .A1(n12), .A2(n141), .ZN(tempResultB[510]) );
  NOR2_X1 U1231 ( .A1(n12), .A2(n144), .ZN(tempResultB[478]) );
  NOR2_X1 U1232 ( .A1(n12), .A2(n147), .ZN(tempResultB[446]) );
  NOR2_X1 U1233 ( .A1(n12), .A2(n150), .ZN(tempResultB[414]) );
  NOR2_X1 U1234 ( .A1(n12), .A2(n153), .ZN(tempResultB[382]) );
  NOR2_X1 U1235 ( .A1(n12), .A2(n156), .ZN(tempResultB[350]) );
  NOR2_X1 U1236 ( .A1(n201), .A2(n186), .ZN(tempResultB[30]) );
  NOR2_X1 U1237 ( .A1(n204), .A2(n189), .ZN(tempResultA_0__26_) );
  NOR2_X1 U1238 ( .A1(n202), .A2(n189), .ZN(tempResultA_0__28_) );
  INV_X1 U1239 ( .A(a_abs[20]), .ZN(n211) );
  NOR2_X1 U1240 ( .A1(n201), .A2(n189), .ZN(tempResultA_0__29_) );
  NOR2_X1 U1241 ( .A1(n210), .A2(n189), .ZN(tempResultA_0__20_) );
  NOR2_X1 U1242 ( .A1(n60), .A2(n140), .ZN(tempResultB[491]) );
  NOR2_X1 U1243 ( .A1(n60), .A2(n143), .ZN(tempResultB[459]) );
  NOR2_X1 U1244 ( .A1(n60), .A2(n146), .ZN(tempResultB[427]) );
  NOR2_X1 U1245 ( .A1(n60), .A2(n149), .ZN(tempResultB[395]) );
  NOR2_X1 U1246 ( .A1(n60), .A2(n152), .ZN(tempResultB[363]) );
  NOR2_X1 U1247 ( .A1(n60), .A2(n155), .ZN(tempResultB[331]) );
  NOR2_X1 U1248 ( .A1(n60), .A2(n185), .ZN(tempResultB[11]) );
  NOR2_X1 U1249 ( .A1(n60), .A2(n188), .ZN(tempResultA_0__10_) );
  NOR2_X1 U1250 ( .A1(n42), .A2(n140), .ZN(tempResultB[497]) );
  NOR2_X1 U1251 ( .A1(n42), .A2(n143), .ZN(tempResultB[465]) );
  NOR2_X1 U1252 ( .A1(n42), .A2(n146), .ZN(tempResultB[433]) );
  NOR2_X1 U1253 ( .A1(n42), .A2(n149), .ZN(tempResultB[401]) );
  NOR2_X1 U1254 ( .A1(n42), .A2(n152), .ZN(tempResultB[369]) );
  NOR2_X1 U1255 ( .A1(n42), .A2(n155), .ZN(tempResultB[337]) );
  NOR2_X1 U1256 ( .A1(n42), .A2(n185), .ZN(tempResultB[17]) );
  NOR2_X1 U1257 ( .A1(n42), .A2(n188), .ZN(tempResultA_0__16_) );
  NOR2_X1 U1258 ( .A1(n20), .A2(n141), .ZN(tempResultB[506]) );
  NOR2_X1 U1259 ( .A1(n20), .A2(n144), .ZN(tempResultB[474]) );
  NOR2_X1 U1260 ( .A1(n20), .A2(n147), .ZN(tempResultB[442]) );
  NOR2_X1 U1261 ( .A1(n20), .A2(n150), .ZN(tempResultB[410]) );
  NOR2_X1 U1262 ( .A1(n20), .A2(n153), .ZN(tempResultB[378]) );
  NOR2_X1 U1263 ( .A1(n20), .A2(n156), .ZN(tempResultB[346]) );
  NOR2_X1 U1264 ( .A1(n205), .A2(n186), .ZN(tempResultB[26]) );
  NOR2_X1 U1265 ( .A1(n205), .A2(n189), .ZN(tempResultA_0__25_) );
  NOR2_X1 U1266 ( .A1(n45), .A2(n140), .ZN(tempResultB[496]) );
  NOR2_X1 U1267 ( .A1(n45), .A2(n143), .ZN(tempResultB[464]) );
  NOR2_X1 U1268 ( .A1(n45), .A2(n146), .ZN(tempResultB[432]) );
  NOR2_X1 U1269 ( .A1(n45), .A2(n149), .ZN(tempResultB[400]) );
  NOR2_X1 U1270 ( .A1(n45), .A2(n152), .ZN(tempResultB[368]) );
  NOR2_X1 U1271 ( .A1(n45), .A2(n155), .ZN(tempResultB[336]) );
  NOR2_X1 U1272 ( .A1(n45), .A2(n185), .ZN(tempResultB[16]) );
  NOR2_X1 U1273 ( .A1(n45), .A2(n188), .ZN(tempResultA_0__15_) );
  NOR2_X1 U1274 ( .A1(n28), .A2(n141), .ZN(tempResultB[502]) );
  NOR2_X1 U1275 ( .A1(n28), .A2(n144), .ZN(tempResultB[470]) );
  NOR2_X1 U1276 ( .A1(n28), .A2(n147), .ZN(tempResultB[438]) );
  NOR2_X1 U1277 ( .A1(n28), .A2(n150), .ZN(tempResultB[406]) );
  NOR2_X1 U1278 ( .A1(n28), .A2(n153), .ZN(tempResultB[374]) );
  NOR2_X1 U1279 ( .A1(n28), .A2(n156), .ZN(tempResultB[342]) );
  NOR2_X1 U1280 ( .A1(n209), .A2(n186), .ZN(tempResultB[22]) );
  NOR2_X1 U1281 ( .A1(n209), .A2(n189), .ZN(tempResultA_0__21_) );
  NOR2_X1 U1282 ( .A1(n22), .A2(n141), .ZN(tempResultB[505]) );
  NOR2_X1 U1283 ( .A1(n22), .A2(n144), .ZN(tempResultB[473]) );
  NOR2_X1 U1284 ( .A1(n22), .A2(n147), .ZN(tempResultB[441]) );
  NOR2_X1 U1285 ( .A1(n22), .A2(n150), .ZN(tempResultB[409]) );
  NOR2_X1 U1286 ( .A1(n22), .A2(n153), .ZN(tempResultB[377]) );
  NOR2_X1 U1287 ( .A1(n22), .A2(n156), .ZN(tempResultB[345]) );
  NOR2_X1 U1288 ( .A1(n206), .A2(n186), .ZN(tempResultB[25]) );
  NOR2_X1 U1289 ( .A1(n24), .A2(n141), .ZN(tempResultB[504]) );
  NOR2_X1 U1290 ( .A1(n24), .A2(n144), .ZN(tempResultB[472]) );
  NOR2_X1 U1291 ( .A1(n24), .A2(n147), .ZN(tempResultB[440]) );
  NOR2_X1 U1292 ( .A1(n24), .A2(n150), .ZN(tempResultB[408]) );
  NOR2_X1 U1293 ( .A1(n24), .A2(n153), .ZN(tempResultB[376]) );
  NOR2_X1 U1294 ( .A1(n24), .A2(n156), .ZN(tempResultB[344]) );
  NOR2_X1 U1295 ( .A1(n207), .A2(n186), .ZN(tempResultB[24]) );
  NOR2_X1 U1296 ( .A1(n207), .A2(n189), .ZN(tempResultA_0__23_) );
  NOR2_X1 U1297 ( .A1(n203), .A2(n189), .ZN(tempResultA_0__27_) );
  NOR2_X1 U1298 ( .A1(n38), .A2(n140), .ZN(tempResultB[498]) );
  NOR2_X1 U1299 ( .A1(n38), .A2(n143), .ZN(tempResultB[466]) );
  NOR2_X1 U1300 ( .A1(n38), .A2(n146), .ZN(tempResultB[434]) );
  NOR2_X1 U1301 ( .A1(n38), .A2(n149), .ZN(tempResultB[402]) );
  NOR2_X1 U1302 ( .A1(n38), .A2(n152), .ZN(tempResultB[370]) );
  NOR2_X1 U1303 ( .A1(n38), .A2(n155), .ZN(tempResultB[338]) );
  NOR2_X1 U1304 ( .A1(n39), .A2(n185), .ZN(tempResultB[18]) );
  NOR2_X1 U1305 ( .A1(n213), .A2(n188), .ZN(tempResultA_0__17_) );
  INV_X1 U1306 ( .A(a_abs[25]), .ZN(n206) );
  NOR2_X1 U1307 ( .A1(n206), .A2(n189), .ZN(tempResultA_0__24_) );
  NOR2_X1 U1308 ( .A1(n66), .A2(n142), .ZN(tempResultB[489]) );
  NOR2_X1 U1309 ( .A1(n66), .A2(n145), .ZN(tempResultB[457]) );
  NOR2_X1 U1310 ( .A1(n66), .A2(n148), .ZN(tempResultB[425]) );
  NOR2_X1 U1311 ( .A1(n66), .A2(n151), .ZN(tempResultB[393]) );
  NOR2_X1 U1312 ( .A1(n66), .A2(n154), .ZN(tempResultB[361]) );
  NOR2_X1 U1313 ( .A1(n66), .A2(n157), .ZN(tempResultB[329]) );
  NOR2_X1 U1314 ( .A1(n66), .A2(n187), .ZN(tempResultB[9]) );
  NOR2_X1 U1315 ( .A1(n66), .A2(n190), .ZN(tempResultA_0__8_) );
  NOR2_X1 U1316 ( .A1(n26), .A2(n141), .ZN(tempResultB[503]) );
  NOR2_X1 U1317 ( .A1(n26), .A2(n144), .ZN(tempResultB[471]) );
  NOR2_X1 U1318 ( .A1(n26), .A2(n147), .ZN(tempResultB[439]) );
  NOR2_X1 U1319 ( .A1(n26), .A2(n150), .ZN(tempResultB[407]) );
  NOR2_X1 U1320 ( .A1(n26), .A2(n153), .ZN(tempResultB[375]) );
  NOR2_X1 U1321 ( .A1(n26), .A2(n156), .ZN(tempResultB[343]) );
  NOR2_X1 U1322 ( .A1(n27), .A2(n186), .ZN(tempResultB[23]) );
  NOR2_X1 U1323 ( .A1(n208), .A2(n189), .ZN(tempResultA_0__22_) );
  NOR2_X1 U1324 ( .A1(n51), .A2(n188), .ZN(tempResultA_0__13_) );
  INV_X1 U1325 ( .A(a_abs[14]), .ZN(n217) );
  INV_X1 U1326 ( .A(a_abs[21]), .ZN(n210) );
  NOR2_X1 U1327 ( .A1(n82), .A2(n142), .ZN(tempResultB[484]) );
  NOR2_X1 U1328 ( .A1(n82), .A2(n145), .ZN(tempResultB[452]) );
  NOR2_X1 U1329 ( .A1(n82), .A2(n148), .ZN(tempResultB[420]) );
  NOR2_X1 U1330 ( .A1(n82), .A2(n151), .ZN(tempResultB[388]) );
  NOR2_X1 U1331 ( .A1(n82), .A2(n154), .ZN(tempResultB[356]) );
  NOR2_X1 U1332 ( .A1(n82), .A2(n157), .ZN(tempResultB[324]) );
  NOR2_X1 U1333 ( .A1(n82), .A2(n187), .ZN(tempResultB[4]) );
  NOR2_X1 U1334 ( .A1(n82), .A2(n190), .ZN(tempResultA_0__3_) );
  NOR2_X1 U1335 ( .A1(n48), .A2(n140), .ZN(tempResultB[495]) );
  NOR2_X1 U1336 ( .A1(n48), .A2(n143), .ZN(tempResultB[463]) );
  NOR2_X1 U1337 ( .A1(n48), .A2(n146), .ZN(tempResultB[431]) );
  NOR2_X1 U1338 ( .A1(n48), .A2(n149), .ZN(tempResultB[399]) );
  NOR2_X1 U1339 ( .A1(n48), .A2(n152), .ZN(tempResultB[367]) );
  NOR2_X1 U1340 ( .A1(n48), .A2(n155), .ZN(tempResultB[335]) );
  NOR2_X1 U1341 ( .A1(n48), .A2(n185), .ZN(tempResultB[15]) );
  NOR2_X1 U1342 ( .A1(n48), .A2(n188), .ZN(tempResultA_0__14_) );
  INV_X1 U1343 ( .A(a_abs[11]), .ZN(n220) );
  NOR2_X1 U1344 ( .A1(n57), .A2(n140), .ZN(tempResultB[492]) );
  NOR2_X1 U1345 ( .A1(n57), .A2(n143), .ZN(tempResultB[460]) );
  NOR2_X1 U1346 ( .A1(n57), .A2(n146), .ZN(tempResultB[428]) );
  NOR2_X1 U1347 ( .A1(n57), .A2(n149), .ZN(tempResultB[396]) );
  NOR2_X1 U1348 ( .A1(n57), .A2(n152), .ZN(tempResultB[364]) );
  NOR2_X1 U1349 ( .A1(n57), .A2(n155), .ZN(tempResultB[332]) );
  NOR2_X1 U1350 ( .A1(n57), .A2(n185), .ZN(tempResultB[12]) );
  NOR2_X1 U1351 ( .A1(n57), .A2(n188), .ZN(tempResultA_0__11_) );
  NOR2_X1 U1352 ( .A1(n70), .A2(n142), .ZN(tempResultB[488]) );
  NOR2_X1 U1353 ( .A1(n70), .A2(n145), .ZN(tempResultB[456]) );
  NOR2_X1 U1354 ( .A1(n70), .A2(n148), .ZN(tempResultB[424]) );
  NOR2_X1 U1355 ( .A1(n70), .A2(n151), .ZN(tempResultB[392]) );
  NOR2_X1 U1356 ( .A1(n70), .A2(n154), .ZN(tempResultB[360]) );
  NOR2_X1 U1357 ( .A1(n70), .A2(n157), .ZN(tempResultB[328]) );
  NOR2_X1 U1358 ( .A1(n70), .A2(n187), .ZN(tempResultB[8]) );
  NOR2_X1 U1359 ( .A1(n70), .A2(n190), .ZN(tempResultA_0__7_) );
  NOR2_X1 U1360 ( .A1(n54), .A2(n140), .ZN(tempResultB[493]) );
  NOR2_X1 U1361 ( .A1(n54), .A2(n143), .ZN(tempResultB[461]) );
  NOR2_X1 U1362 ( .A1(n54), .A2(n146), .ZN(tempResultB[429]) );
  NOR2_X1 U1363 ( .A1(n54), .A2(n149), .ZN(tempResultB[397]) );
  NOR2_X1 U1364 ( .A1(n54), .A2(n152), .ZN(tempResultB[365]) );
  NOR2_X1 U1365 ( .A1(n54), .A2(n155), .ZN(tempResultB[333]) );
  NOR2_X1 U1366 ( .A1(n54), .A2(n185), .ZN(tempResultB[13]) );
  NOR2_X1 U1367 ( .A1(n54), .A2(n188), .ZN(tempResultA_0__12_) );
  NOR2_X1 U1368 ( .A1(n73), .A2(n142), .ZN(tempResultB[487]) );
  NOR2_X1 U1369 ( .A1(n73), .A2(n145), .ZN(tempResultB[455]) );
  NOR2_X1 U1370 ( .A1(n73), .A2(n148), .ZN(tempResultB[423]) );
  NOR2_X1 U1371 ( .A1(n73), .A2(n151), .ZN(tempResultB[391]) );
  NOR2_X1 U1372 ( .A1(n73), .A2(n154), .ZN(tempResultB[359]) );
  NOR2_X1 U1373 ( .A1(n73), .A2(n157), .ZN(tempResultB[327]) );
  NOR2_X1 U1374 ( .A1(n73), .A2(n187), .ZN(tempResultB[7]) );
  NOR2_X1 U1375 ( .A1(n73), .A2(n190), .ZN(tempResultA_0__6_) );
  INV_X1 U1376 ( .A(a_abs[9]), .ZN(n222) );
  NOR2_X1 U1377 ( .A1(n79), .A2(n142), .ZN(tempResultB[485]) );
  NOR2_X1 U1378 ( .A1(n79), .A2(n145), .ZN(tempResultB[453]) );
  NOR2_X1 U1379 ( .A1(n79), .A2(n148), .ZN(tempResultB[421]) );
  NOR2_X1 U1380 ( .A1(n79), .A2(n151), .ZN(tempResultB[389]) );
  NOR2_X1 U1381 ( .A1(n79), .A2(n154), .ZN(tempResultB[357]) );
  NOR2_X1 U1382 ( .A1(n79), .A2(n157), .ZN(tempResultB[325]) );
  NOR2_X1 U1383 ( .A1(n79), .A2(n187), .ZN(tempResultB[5]) );
  NOR2_X1 U1384 ( .A1(n79), .A2(n190), .ZN(tempResultA_0__4_) );
  NOR2_X1 U1385 ( .A1(n76), .A2(n142), .ZN(tempResultB[486]) );
  NOR2_X1 U1386 ( .A1(n76), .A2(n145), .ZN(tempResultB[454]) );
  NOR2_X1 U1387 ( .A1(n76), .A2(n148), .ZN(tempResultB[422]) );
  NOR2_X1 U1388 ( .A1(n76), .A2(n151), .ZN(tempResultB[390]) );
  NOR2_X1 U1389 ( .A1(n76), .A2(n154), .ZN(tempResultB[358]) );
  NOR2_X1 U1390 ( .A1(n76), .A2(n157), .ZN(tempResultB[326]) );
  NOR2_X1 U1391 ( .A1(n76), .A2(n187), .ZN(tempResultB[6]) );
  NOR2_X1 U1392 ( .A1(n76), .A2(n190), .ZN(tempResultA_0__5_) );
  INV_X1 U1393 ( .A(a_abs[7]), .ZN(n224) );
  INV_X1 U1394 ( .A(a_abs[4]), .ZN(n227) );
  NOR2_X1 U1395 ( .A1(n85), .A2(n142), .ZN(tempResultB[483]) );
  NOR2_X1 U1396 ( .A1(n85), .A2(n145), .ZN(tempResultB[451]) );
  NOR2_X1 U1397 ( .A1(n85), .A2(n148), .ZN(tempResultB[419]) );
  NOR2_X1 U1398 ( .A1(n85), .A2(n151), .ZN(tempResultB[387]) );
  NOR2_X1 U1399 ( .A1(n85), .A2(n154), .ZN(tempResultB[355]) );
  NOR2_X1 U1400 ( .A1(n85), .A2(n157), .ZN(tempResultB[323]) );
  NOR2_X1 U1401 ( .A1(n85), .A2(n187), .ZN(tempResultB[3]) );
  NOR2_X1 U1402 ( .A1(n85), .A2(n189), .ZN(tempResultA_0__2_) );
  NOR2_X1 U1403 ( .A1(n88), .A2(n141), .ZN(tempResultB[482]) );
  NOR2_X1 U1404 ( .A1(n88), .A2(n144), .ZN(tempResultB[450]) );
  NOR2_X1 U1405 ( .A1(n88), .A2(n147), .ZN(tempResultB[418]) );
  NOR2_X1 U1406 ( .A1(n88), .A2(n150), .ZN(tempResultB[386]) );
  NOR2_X1 U1407 ( .A1(n88), .A2(n153), .ZN(tempResultB[354]) );
  NOR2_X1 U1408 ( .A1(n88), .A2(n156), .ZN(tempResultB[322]) );
  NOR2_X1 U1409 ( .A1(n88), .A2(n186), .ZN(tempResultB[2]) );
  NOR2_X1 U1410 ( .A1(n88), .A2(n189), .ZN(tempResultA_0__1_) );
  BUF_X4 U1411 ( .A(b[31]), .Z(n197) );
  BUF_X4 U1412 ( .A(b[31]), .Z(n198) );
  BUF_X1 U1413 ( .A(finalSign), .Z(n191) );
  BUF_X1 U1414 ( .A(finalSign), .Z(n192) );
endmodule


module register_N64 ( clk, reset, reg_in, reg_out );
  input [63:0] reg_in;
  output [63:0] reg_out;
  input clk, reset;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73;

  SDFF_X1 reg_out_reg_63_ ( .D(1'b0), .SI(n65), .SE(reg_in[63]), .CK(clk), .Q(
        reg_out[63]) );
  SDFF_X1 reg_out_reg_62_ ( .D(1'b0), .SI(n65), .SE(reg_in[62]), .CK(clk), .Q(
        reg_out[62]) );
  SDFF_X1 reg_out_reg_61_ ( .D(1'b0), .SI(n65), .SE(reg_in[61]), .CK(clk), .Q(
        reg_out[61]) );
  SDFF_X1 reg_out_reg_60_ ( .D(1'b0), .SI(n65), .SE(reg_in[60]), .CK(clk), .Q(
        reg_out[60]) );
  SDFF_X1 reg_out_reg_59_ ( .D(1'b0), .SI(n65), .SE(reg_in[59]), .CK(clk), .Q(
        reg_out[59]) );
  SDFF_X1 reg_out_reg_58_ ( .D(1'b0), .SI(n65), .SE(reg_in[58]), .CK(clk), .Q(
        reg_out[58]) );
  SDFF_X1 reg_out_reg_57_ ( .D(1'b0), .SI(n65), .SE(reg_in[57]), .CK(clk), .Q(
        reg_out[57]) );
  SDFF_X1 reg_out_reg_56_ ( .D(1'b0), .SI(n65), .SE(reg_in[56]), .CK(clk), .Q(
        reg_out[56]) );
  SDFF_X1 reg_out_reg_55_ ( .D(1'b0), .SI(n65), .SE(reg_in[55]), .CK(clk), .Q(
        reg_out[55]) );
  SDFF_X1 reg_out_reg_54_ ( .D(1'b0), .SI(n65), .SE(reg_in[54]), .CK(clk), .Q(
        reg_out[54]) );
  SDFF_X1 reg_out_reg_53_ ( .D(1'b0), .SI(n65), .SE(reg_in[53]), .CK(clk), .Q(
        reg_out[53]) );
  SDFF_X1 reg_out_reg_52_ ( .D(1'b0), .SI(n66), .SE(reg_in[52]), .CK(clk), .Q(
        reg_out[52]) );
  SDFF_X1 reg_out_reg_51_ ( .D(1'b0), .SI(n66), .SE(reg_in[51]), .CK(clk), .Q(
        reg_out[51]) );
  SDFF_X1 reg_out_reg_50_ ( .D(1'b0), .SI(n66), .SE(reg_in[50]), .CK(clk), .Q(
        reg_out[50]) );
  SDFF_X1 reg_out_reg_49_ ( .D(1'b0), .SI(n66), .SE(reg_in[49]), .CK(clk), .Q(
        reg_out[49]) );
  SDFF_X1 reg_out_reg_48_ ( .D(1'b0), .SI(n66), .SE(reg_in[48]), .CK(clk), .Q(
        reg_out[48]) );
  SDFF_X1 reg_out_reg_47_ ( .D(1'b0), .SI(n66), .SE(reg_in[47]), .CK(clk), .Q(
        reg_out[47]) );
  SDFF_X1 reg_out_reg_46_ ( .D(1'b0), .SI(n66), .SE(reg_in[46]), .CK(clk), .Q(
        reg_out[46]) );
  SDFF_X1 reg_out_reg_45_ ( .D(1'b0), .SI(n66), .SE(reg_in[45]), .CK(clk), .Q(
        reg_out[45]) );
  SDFF_X1 reg_out_reg_44_ ( .D(1'b0), .SI(n66), .SE(reg_in[44]), .CK(clk), .Q(
        reg_out[44]) );
  SDFF_X1 reg_out_reg_43_ ( .D(1'b0), .SI(n66), .SE(reg_in[43]), .CK(clk), .Q(
        reg_out[43]) );
  SDFF_X1 reg_out_reg_42_ ( .D(1'b0), .SI(n66), .SE(reg_in[42]), .CK(clk), .Q(
        reg_out[42]) );
  SDFF_X1 reg_out_reg_41_ ( .D(1'b0), .SI(n67), .SE(reg_in[41]), .CK(clk), .Q(
        reg_out[41]) );
  SDFF_X1 reg_out_reg_40_ ( .D(1'b0), .SI(n67), .SE(reg_in[40]), .CK(clk), .Q(
        reg_out[40]) );
  SDFF_X1 reg_out_reg_39_ ( .D(1'b0), .SI(n67), .SE(reg_in[39]), .CK(clk), .Q(
        reg_out[39]) );
  SDFF_X1 reg_out_reg_38_ ( .D(1'b0), .SI(n67), .SE(reg_in[38]), .CK(clk), .Q(
        reg_out[38]) );
  SDFF_X1 reg_out_reg_37_ ( .D(1'b0), .SI(n67), .SE(reg_in[37]), .CK(clk), .Q(
        reg_out[37]) );
  SDFF_X1 reg_out_reg_36_ ( .D(1'b0), .SI(n67), .SE(reg_in[36]), .CK(clk), .Q(
        reg_out[36]) );
  SDFF_X1 reg_out_reg_35_ ( .D(1'b0), .SI(n67), .SE(reg_in[35]), .CK(clk), .Q(
        reg_out[35]) );
  SDFF_X1 reg_out_reg_34_ ( .D(1'b0), .SI(n67), .SE(reg_in[34]), .CK(clk), .Q(
        reg_out[34]) );
  SDFF_X1 reg_out_reg_33_ ( .D(1'b0), .SI(n67), .SE(reg_in[33]), .CK(clk), .Q(
        reg_out[33]) );
  SDFF_X1 reg_out_reg_32_ ( .D(1'b0), .SI(n67), .SE(reg_in[32]), .CK(clk), .Q(
        reg_out[32]) );
  SDFF_X1 reg_out_reg_31_ ( .D(1'b0), .SI(n67), .SE(reg_in[31]), .CK(clk), .Q(
        reg_out[31]) );
  SDFF_X1 reg_out_reg_30_ ( .D(1'b0), .SI(n68), .SE(reg_in[30]), .CK(clk), .Q(
        reg_out[30]) );
  SDFF_X1 reg_out_reg_29_ ( .D(1'b0), .SI(n68), .SE(reg_in[29]), .CK(clk), .Q(
        reg_out[29]) );
  SDFF_X1 reg_out_reg_28_ ( .D(1'b0), .SI(n68), .SE(reg_in[28]), .CK(clk), .Q(
        reg_out[28]) );
  SDFF_X1 reg_out_reg_27_ ( .D(1'b0), .SI(n68), .SE(reg_in[27]), .CK(clk), .Q(
        reg_out[27]) );
  SDFF_X1 reg_out_reg_26_ ( .D(1'b0), .SI(n68), .SE(reg_in[26]), .CK(clk), .Q(
        reg_out[26]) );
  SDFF_X1 reg_out_reg_25_ ( .D(1'b0), .SI(n68), .SE(reg_in[25]), .CK(clk), .Q(
        reg_out[25]) );
  SDFF_X1 reg_out_reg_24_ ( .D(1'b0), .SI(n68), .SE(reg_in[24]), .CK(clk), .Q(
        reg_out[24]) );
  SDFF_X1 reg_out_reg_23_ ( .D(1'b0), .SI(n68), .SE(reg_in[23]), .CK(clk), .Q(
        reg_out[23]) );
  SDFF_X1 reg_out_reg_22_ ( .D(1'b0), .SI(n68), .SE(reg_in[22]), .CK(clk), .Q(
        reg_out[22]) );
  SDFF_X1 reg_out_reg_21_ ( .D(1'b0), .SI(n68), .SE(reg_in[21]), .CK(clk), .Q(
        reg_out[21]) );
  SDFF_X1 reg_out_reg_20_ ( .D(1'b0), .SI(n68), .SE(reg_in[20]), .CK(clk), .Q(
        reg_out[20]) );
  SDFF_X1 reg_out_reg_19_ ( .D(1'b0), .SI(n69), .SE(reg_in[19]), .CK(clk), .Q(
        reg_out[19]) );
  SDFF_X1 reg_out_reg_18_ ( .D(1'b0), .SI(n69), .SE(reg_in[18]), .CK(clk), .Q(
        reg_out[18]) );
  SDFF_X1 reg_out_reg_17_ ( .D(1'b0), .SI(n69), .SE(reg_in[17]), .CK(clk), .Q(
        reg_out[17]) );
  SDFF_X1 reg_out_reg_16_ ( .D(1'b0), .SI(n69), .SE(reg_in[16]), .CK(clk), .Q(
        reg_out[16]) );
  SDFF_X1 reg_out_reg_15_ ( .D(1'b0), .SI(n69), .SE(reg_in[15]), .CK(clk), .Q(
        reg_out[15]) );
  SDFF_X1 reg_out_reg_14_ ( .D(1'b0), .SI(n69), .SE(reg_in[14]), .CK(clk), .Q(
        reg_out[14]) );
  SDFF_X1 reg_out_reg_13_ ( .D(1'b0), .SI(n69), .SE(reg_in[13]), .CK(clk), .Q(
        reg_out[13]) );
  SDFF_X1 reg_out_reg_12_ ( .D(1'b0), .SI(n69), .SE(reg_in[12]), .CK(clk), .Q(
        reg_out[12]) );
  SDFF_X1 reg_out_reg_11_ ( .D(1'b0), .SI(n69), .SE(reg_in[11]), .CK(clk), .Q(
        reg_out[11]) );
  SDFF_X1 reg_out_reg_10_ ( .D(1'b0), .SI(n69), .SE(reg_in[10]), .CK(clk), .Q(
        reg_out[10]) );
  SDFF_X1 reg_out_reg_9_ ( .D(1'b0), .SI(n69), .SE(reg_in[9]), .CK(clk), .Q(
        reg_out[9]) );
  SDFF_X1 reg_out_reg_8_ ( .D(1'b0), .SI(n70), .SE(reg_in[8]), .CK(clk), .Q(
        reg_out[8]) );
  SDFF_X1 reg_out_reg_7_ ( .D(1'b0), .SI(n70), .SE(reg_in[7]), .CK(clk), .Q(
        reg_out[7]) );
  SDFF_X1 reg_out_reg_6_ ( .D(1'b0), .SI(n70), .SE(reg_in[6]), .CK(clk), .Q(
        reg_out[6]) );
  SDFF_X1 reg_out_reg_5_ ( .D(1'b0), .SI(n70), .SE(reg_in[5]), .CK(clk), .Q(
        reg_out[5]) );
  SDFF_X1 reg_out_reg_4_ ( .D(1'b0), .SI(n70), .SE(reg_in[4]), .CK(clk), .Q(
        reg_out[4]) );
  SDFF_X1 reg_out_reg_3_ ( .D(1'b0), .SI(n70), .SE(reg_in[3]), .CK(clk), .Q(
        reg_out[3]) );
  SDFF_X1 reg_out_reg_2_ ( .D(1'b0), .SI(n70), .SE(reg_in[2]), .CK(clk), .Q(
        reg_out[2]) );
  SDFF_X1 reg_out_reg_1_ ( .D(1'b0), .SI(n70), .SE(reg_in[1]), .CK(clk), .Q(
        reg_out[1]) );
  SDFF_X1 reg_out_reg_0_ ( .D(1'b0), .SI(n70), .SE(reg_in[0]), .CK(clk), .Q(
        reg_out[0]) );
  BUF_X1 U67 ( .A(n71), .Z(n69) );
  BUF_X1 U68 ( .A(n71), .Z(n68) );
  BUF_X1 U69 ( .A(n72), .Z(n67) );
  BUF_X1 U70 ( .A(n72), .Z(n66) );
  BUF_X1 U71 ( .A(n72), .Z(n65) );
  BUF_X1 U72 ( .A(n71), .Z(n70) );
  INV_X1 U73 ( .A(reset), .ZN(n73) );
  BUF_X1 U74 ( .A(n73), .Z(n71) );
  BUF_X1 U75 ( .A(n73), .Z(n72) );
endmodule


module TopModule ( clk, a, b, reset, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;
  input clk, reset;

  wire   [31:0] mulA;
  wire   [31:0] mulB;
  wire   [63:0] mulResult;

  register_N32_0 R0 ( .clk(clk), .reset(reset), .reg_in(a), .reg_out(mulA) );
  register_N32_1 R1 ( .clk(clk), .reset(reset), .reg_in(b), .reg_out(mulB) );
  multiplierTreeV2 M0 ( .a(mulA), .b(mulB), .result(mulResult) );
  register_N64 R2 ( .clk(clk), .reset(reset), .reg_in(mulResult), .reg_out(
        result) );
endmodule

